module STORE_QUEUE_LSQ_dist( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_bbStart, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_0, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_1, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_2, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_3, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_4, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_5, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_6, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_7, // @[:@6.4]
  input  [2:0]  io_bbNumStores, // @[:@6.4]
  output [2:0]  io_storeTail, // @[:@6.4]
  output [2:0]  io_storeHead, // @[:@6.4]
  output        io_storeEmpty, // @[:@6.4]
  input  [2:0]  io_loadTail, // @[:@6.4]
  input  [2:0]  io_loadHead, // @[:@6.4]
  input         io_loadEmpty, // @[:@6.4]
  input         io_loadAddressDone_0, // @[:@6.4]
  input         io_loadAddressDone_1, // @[:@6.4]
  input         io_loadAddressDone_2, // @[:@6.4]
  input         io_loadAddressDone_3, // @[:@6.4]
  input         io_loadAddressDone_4, // @[:@6.4]
  input         io_loadAddressDone_5, // @[:@6.4]
  input         io_loadAddressDone_6, // @[:@6.4]
  input         io_loadAddressDone_7, // @[:@6.4]
  input         io_loadDataDone_0, // @[:@6.4]
  input         io_loadDataDone_1, // @[:@6.4]
  input         io_loadDataDone_2, // @[:@6.4]
  input         io_loadDataDone_3, // @[:@6.4]
  input         io_loadDataDone_4, // @[:@6.4]
  input         io_loadDataDone_5, // @[:@6.4]
  input         io_loadDataDone_6, // @[:@6.4]
  input         io_loadDataDone_7, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_0, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_1, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_2, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_3, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_4, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_5, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_6, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_7, // @[:@6.4]
  output        io_storeAddrDone_0, // @[:@6.4]
  output        io_storeAddrDone_1, // @[:@6.4]
  output        io_storeAddrDone_2, // @[:@6.4]
  output        io_storeAddrDone_3, // @[:@6.4]
  output        io_storeAddrDone_4, // @[:@6.4]
  output        io_storeAddrDone_5, // @[:@6.4]
  output        io_storeAddrDone_6, // @[:@6.4]
  output        io_storeAddrDone_7, // @[:@6.4]
  output        io_storeDataDone_0, // @[:@6.4]
  output        io_storeDataDone_1, // @[:@6.4]
  output        io_storeDataDone_2, // @[:@6.4]
  output        io_storeDataDone_3, // @[:@6.4]
  output        io_storeDataDone_4, // @[:@6.4]
  output        io_storeDataDone_5, // @[:@6.4]
  output        io_storeDataDone_6, // @[:@6.4]
  output        io_storeDataDone_7, // @[:@6.4]
  output [31:0] io_storeAddrQueue_0, // @[:@6.4]
  output [31:0] io_storeAddrQueue_1, // @[:@6.4]
  output [31:0] io_storeAddrQueue_2, // @[:@6.4]
  output [31:0] io_storeAddrQueue_3, // @[:@6.4]
  output [31:0] io_storeAddrQueue_4, // @[:@6.4]
  output [31:0] io_storeAddrQueue_5, // @[:@6.4]
  output [31:0] io_storeAddrQueue_6, // @[:@6.4]
  output [31:0] io_storeAddrQueue_7, // @[:@6.4]
  output [31:0] io_storeDataQueue_0, // @[:@6.4]
  output [31:0] io_storeDataQueue_1, // @[:@6.4]
  output [31:0] io_storeDataQueue_2, // @[:@6.4]
  output [31:0] io_storeDataQueue_3, // @[:@6.4]
  output [31:0] io_storeDataQueue_4, // @[:@6.4]
  output [31:0] io_storeDataQueue_5, // @[:@6.4]
  output [31:0] io_storeDataQueue_6, // @[:@6.4]
  output [31:0] io_storeDataQueue_7, // @[:@6.4]
  input         io_storeDataEnable_0, // @[:@6.4]
  input  [31:0] io_dataFromStorePorts_0, // @[:@6.4]
  input         io_storeAddrEnable_0, // @[:@6.4]
  input  [31:0] io_addressFromStorePorts_0, // @[:@6.4]
  output [31:0] io_storeAddrToMem, // @[:@6.4]
  output [31:0] io_storeDataToMem, // @[:@6.4]
  output        io_storeEnableToMem, // @[:@6.4]
  input         io_memIsReadyForStores // @[:@6.4]
);
  reg [2:0] head; // @[StoreQueue.scala 50:21:@8.4]
  reg [31:0] _RAND_0;
  reg [2:0] tail; // @[StoreQueue.scala 51:21:@9.4]
  reg [31:0] _RAND_1;
  reg [2:0] offsetQ_0; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_2;
  reg [2:0] offsetQ_1; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_3;
  reg [2:0] offsetQ_2; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_4;
  reg [2:0] offsetQ_3; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_5;
  reg [2:0] offsetQ_4; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_6;
  reg [2:0] offsetQ_5; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_7;
  reg [2:0] offsetQ_6; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_8;
  reg [2:0] offsetQ_7; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_9;
  reg  portQ_0; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_10;
  reg  portQ_1; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_11;
  reg  portQ_2; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_12;
  reg  portQ_3; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_13;
  reg  portQ_4; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_14;
  reg  portQ_5; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_15;
  reg  portQ_6; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_16;
  reg  portQ_7; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_17;
  reg [31:0] addrQ_0; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_18;
  reg [31:0] addrQ_1; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_19;
  reg [31:0] addrQ_2; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_20;
  reg [31:0] addrQ_3; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_21;
  reg [31:0] addrQ_4; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_22;
  reg [31:0] addrQ_5; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_23;
  reg [31:0] addrQ_6; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_24;
  reg [31:0] addrQ_7; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_25;
  reg [31:0] dataQ_0; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_26;
  reg [31:0] dataQ_1; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_27;
  reg [31:0] dataQ_2; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_28;
  reg [31:0] dataQ_3; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_29;
  reg [31:0] dataQ_4; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_30;
  reg [31:0] dataQ_5; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_31;
  reg [31:0] dataQ_6; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_32;
  reg [31:0] dataQ_7; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_33;
  reg  addrKnown_0; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_34;
  reg  addrKnown_1; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_35;
  reg  addrKnown_2; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_36;
  reg  addrKnown_3; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_37;
  reg  addrKnown_4; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_38;
  reg  addrKnown_5; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_39;
  reg  addrKnown_6; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_40;
  reg  addrKnown_7; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_41;
  reg  dataKnown_0; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_42;
  reg  dataKnown_1; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_43;
  reg  dataKnown_2; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_44;
  reg  dataKnown_3; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_45;
  reg  dataKnown_4; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_46;
  reg  dataKnown_5; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_47;
  reg  dataKnown_6; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_48;
  reg  dataKnown_7; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_49;
  reg  allocatedEntries_0; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_50;
  reg  allocatedEntries_1; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_51;
  reg  allocatedEntries_2; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_52;
  reg  allocatedEntries_3; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_53;
  reg  allocatedEntries_4; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_54;
  reg  allocatedEntries_5; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_55;
  reg  allocatedEntries_6; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_56;
  reg  allocatedEntries_7; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_57;
  reg  storeCompleted_0; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_58;
  reg  storeCompleted_1; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_59;
  reg  storeCompleted_2; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_60;
  reg  storeCompleted_3; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_61;
  reg  storeCompleted_4; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_62;
  reg  storeCompleted_5; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_63;
  reg  storeCompleted_6; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_64;
  reg  storeCompleted_7; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_65;
  reg  checkBits_0; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_66;
  reg  checkBits_1; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_67;
  reg  checkBits_2; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_68;
  reg  checkBits_3; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_69;
  reg  checkBits_4; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_70;
  reg  checkBits_5; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_71;
  reg  checkBits_6; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_72;
  reg  checkBits_7; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_73;
  wire [4:0] _GEN_378; // @[util.scala 14:20:@101.4]
  wire [5:0] _T_948; // @[util.scala 14:20:@101.4]
  wire [5:0] _T_949; // @[util.scala 14:20:@102.4]
  wire [4:0] _T_950; // @[util.scala 14:20:@103.4]
  wire [4:0] _GEN_0; // @[util.scala 14:25:@104.4]
  wire [3:0] _T_951; // @[util.scala 14:25:@104.4]
  wire [3:0] _GEN_379; // @[StoreQueue.scala 70:46:@105.4]
  wire  _T_952; // @[StoreQueue.scala 70:46:@105.4]
  wire  initBits_0; // @[StoreQueue.scala 70:64:@106.4]
  wire [5:0] _T_957; // @[util.scala 14:20:@108.4]
  wire [5:0] _T_958; // @[util.scala 14:20:@109.4]
  wire [4:0] _T_959; // @[util.scala 14:20:@110.4]
  wire [4:0] _GEN_8; // @[util.scala 14:25:@111.4]
  wire [3:0] _T_960; // @[util.scala 14:25:@111.4]
  wire  _T_961; // @[StoreQueue.scala 70:46:@112.4]
  wire  initBits_1; // @[StoreQueue.scala 70:64:@113.4]
  wire [5:0] _T_966; // @[util.scala 14:20:@115.4]
  wire [5:0] _T_967; // @[util.scala 14:20:@116.4]
  wire [4:0] _T_968; // @[util.scala 14:20:@117.4]
  wire [4:0] _GEN_9; // @[util.scala 14:25:@118.4]
  wire [3:0] _T_969; // @[util.scala 14:25:@118.4]
  wire  _T_970; // @[StoreQueue.scala 70:46:@119.4]
  wire  initBits_2; // @[StoreQueue.scala 70:64:@120.4]
  wire [5:0] _T_975; // @[util.scala 14:20:@122.4]
  wire [5:0] _T_976; // @[util.scala 14:20:@123.4]
  wire [4:0] _T_977; // @[util.scala 14:20:@124.4]
  wire [4:0] _GEN_10; // @[util.scala 14:25:@125.4]
  wire [3:0] _T_978; // @[util.scala 14:25:@125.4]
  wire  _T_979; // @[StoreQueue.scala 70:46:@126.4]
  wire  initBits_3; // @[StoreQueue.scala 70:64:@127.4]
  wire [5:0] _T_984; // @[util.scala 14:20:@129.4]
  wire [5:0] _T_985; // @[util.scala 14:20:@130.4]
  wire [4:0] _T_986; // @[util.scala 14:20:@131.4]
  wire [4:0] _GEN_11; // @[util.scala 14:25:@132.4]
  wire [3:0] _T_987; // @[util.scala 14:25:@132.4]
  wire  _T_988; // @[StoreQueue.scala 70:46:@133.4]
  wire  initBits_4; // @[StoreQueue.scala 70:64:@134.4]
  wire [5:0] _T_993; // @[util.scala 14:20:@136.4]
  wire [5:0] _T_994; // @[util.scala 14:20:@137.4]
  wire [4:0] _T_995; // @[util.scala 14:20:@138.4]
  wire [4:0] _GEN_12; // @[util.scala 14:25:@139.4]
  wire [3:0] _T_996; // @[util.scala 14:25:@139.4]
  wire  _T_997; // @[StoreQueue.scala 70:46:@140.4]
  wire  initBits_5; // @[StoreQueue.scala 70:64:@141.4]
  wire [5:0] _T_1002; // @[util.scala 14:20:@143.4]
  wire [5:0] _T_1003; // @[util.scala 14:20:@144.4]
  wire [4:0] _T_1004; // @[util.scala 14:20:@145.4]
  wire [4:0] _GEN_13; // @[util.scala 14:25:@146.4]
  wire [3:0] _T_1005; // @[util.scala 14:25:@146.4]
  wire  _T_1006; // @[StoreQueue.scala 70:46:@147.4]
  wire  initBits_6; // @[StoreQueue.scala 70:64:@148.4]
  wire [5:0] _T_1011; // @[util.scala 14:20:@150.4]
  wire [5:0] _T_1012; // @[util.scala 14:20:@151.4]
  wire [4:0] _T_1013; // @[util.scala 14:20:@152.4]
  wire [4:0] _GEN_14; // @[util.scala 14:25:@153.4]
  wire [3:0] _T_1014; // @[util.scala 14:25:@153.4]
  wire  _T_1015; // @[StoreQueue.scala 70:46:@154.4]
  wire  initBits_7; // @[StoreQueue.scala 70:64:@155.4]
  wire  _T_1030; // @[StoreQueue.scala 72:78:@165.4]
  wire  _T_1031; // @[StoreQueue.scala 72:78:@166.4]
  wire  _T_1032; // @[StoreQueue.scala 72:78:@167.4]
  wire  _T_1033; // @[StoreQueue.scala 72:78:@168.4]
  wire  _T_1034; // @[StoreQueue.scala 72:78:@169.4]
  wire  _T_1035; // @[StoreQueue.scala 72:78:@170.4]
  wire  _T_1036; // @[StoreQueue.scala 72:78:@171.4]
  wire  _T_1037; // @[StoreQueue.scala 72:78:@172.4]
  wire [2:0] _T_1060; // @[:@196.6]
  wire [2:0] _GEN_1; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_2; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_3; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_4; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_5; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_6; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_7; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_16; // @[StoreQueue.scala 75:25:@190.4]
  wire  _GEN_17; // @[StoreQueue.scala 75:25:@190.4]
  wire [2:0] _T_1078; // @[:@212.6]
  wire [2:0] _GEN_19; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_20; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_21; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_22; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_23; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_24; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_25; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_34; // @[StoreQueue.scala 75:25:@206.4]
  wire  _GEN_35; // @[StoreQueue.scala 75:25:@206.4]
  wire [2:0] _T_1096; // @[:@228.6]
  wire [2:0] _GEN_37; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_38; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_39; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_40; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_41; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_42; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_43; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_52; // @[StoreQueue.scala 75:25:@222.4]
  wire  _GEN_53; // @[StoreQueue.scala 75:25:@222.4]
  wire [2:0] _T_1114; // @[:@244.6]
  wire [2:0] _GEN_55; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_56; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_57; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_58; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_59; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_60; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_61; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_70; // @[StoreQueue.scala 75:25:@238.4]
  wire  _GEN_71; // @[StoreQueue.scala 75:25:@238.4]
  wire [2:0] _T_1132; // @[:@260.6]
  wire [2:0] _GEN_73; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_74; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_75; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_76; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_77; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_78; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_79; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_88; // @[StoreQueue.scala 75:25:@254.4]
  wire  _GEN_89; // @[StoreQueue.scala 75:25:@254.4]
  wire [2:0] _T_1150; // @[:@276.6]
  wire [2:0] _GEN_91; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_92; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_93; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_94; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_95; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_96; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_97; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_106; // @[StoreQueue.scala 75:25:@270.4]
  wire  _GEN_107; // @[StoreQueue.scala 75:25:@270.4]
  wire [2:0] _T_1168; // @[:@292.6]
  wire [2:0] _GEN_109; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_110; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_111; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_112; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_113; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_114; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_115; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_124; // @[StoreQueue.scala 75:25:@286.4]
  wire  _GEN_125; // @[StoreQueue.scala 75:25:@286.4]
  wire [2:0] _T_1186; // @[:@308.6]
  wire [2:0] _GEN_127; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_128; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_129; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_130; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_131; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_132; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_133; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_142; // @[StoreQueue.scala 75:25:@302.4]
  wire  _GEN_143; // @[StoreQueue.scala 75:25:@302.4]
  reg [2:0] previousLoadHead; // @[StoreQueue.scala 92:33:@318.4]
  reg [31:0] _RAND_74;
  wire [3:0] _T_1208; // @[util.scala 10:8:@327.6]
  wire [3:0] _GEN_15; // @[util.scala 10:14:@328.6]
  wire [3:0] _T_1209; // @[util.scala 10:14:@328.6]
  wire [3:0] _GEN_411; // @[StoreQueue.scala 96:56:@329.6]
  wire  _T_1210; // @[StoreQueue.scala 96:56:@329.6]
  wire  _T_1211; // @[StoreQueue.scala 95:50:@330.6]
  wire  _T_1213; // @[StoreQueue.scala 95:35:@331.6]
  wire  _T_1215; // @[StoreQueue.scala 100:35:@339.8]
  wire  _T_1216; // @[StoreQueue.scala 100:87:@340.8]
  wire  _T_1217; // @[StoreQueue.scala 100:61:@341.8]
  wire  _T_1219; // @[StoreQueue.scala 102:35:@346.10]
  wire  _T_1220; // @[StoreQueue.scala 103:23:@347.10]
  wire  _T_1221; // @[StoreQueue.scala 103:75:@348.10]
  wire  _T_1222; // @[StoreQueue.scala 103:49:@349.10]
  wire  _T_1224; // @[StoreQueue.scala 103:9:@350.10]
  wire  _T_1225; // @[StoreQueue.scala 102:49:@351.10]
  wire  _GEN_152; // @[StoreQueue.scala 103:96:@352.10]
  wire  _GEN_153; // @[StoreQueue.scala 100:102:@342.8]
  wire  _GEN_154; // @[StoreQueue.scala 98:26:@335.6]
  wire  _GEN_155; // @[StoreQueue.scala 94:35:@320.4]
  wire [3:0] _T_1238; // @[util.scala 10:8:@363.6]
  wire [3:0] _GEN_18; // @[util.scala 10:14:@364.6]
  wire [3:0] _T_1239; // @[util.scala 10:14:@364.6]
  wire  _T_1240; // @[StoreQueue.scala 96:56:@365.6]
  wire  _T_1241; // @[StoreQueue.scala 95:50:@366.6]
  wire  _T_1243; // @[StoreQueue.scala 95:35:@367.6]
  wire  _T_1245; // @[StoreQueue.scala 100:35:@375.8]
  wire  _T_1246; // @[StoreQueue.scala 100:87:@376.8]
  wire  _T_1247; // @[StoreQueue.scala 100:61:@377.8]
  wire  _T_1250; // @[StoreQueue.scala 103:23:@383.10]
  wire  _T_1251; // @[StoreQueue.scala 103:75:@384.10]
  wire  _T_1252; // @[StoreQueue.scala 103:49:@385.10]
  wire  _T_1254; // @[StoreQueue.scala 103:9:@386.10]
  wire  _T_1255; // @[StoreQueue.scala 102:49:@387.10]
  wire  _GEN_164; // @[StoreQueue.scala 103:96:@388.10]
  wire  _GEN_165; // @[StoreQueue.scala 100:102:@378.8]
  wire  _GEN_166; // @[StoreQueue.scala 98:26:@371.6]
  wire  _GEN_167; // @[StoreQueue.scala 94:35:@356.4]
  wire [3:0] _T_1268; // @[util.scala 10:8:@399.6]
  wire [3:0] _GEN_26; // @[util.scala 10:14:@400.6]
  wire [3:0] _T_1269; // @[util.scala 10:14:@400.6]
  wire  _T_1270; // @[StoreQueue.scala 96:56:@401.6]
  wire  _T_1271; // @[StoreQueue.scala 95:50:@402.6]
  wire  _T_1273; // @[StoreQueue.scala 95:35:@403.6]
  wire  _T_1275; // @[StoreQueue.scala 100:35:@411.8]
  wire  _T_1276; // @[StoreQueue.scala 100:87:@412.8]
  wire  _T_1277; // @[StoreQueue.scala 100:61:@413.8]
  wire  _T_1280; // @[StoreQueue.scala 103:23:@419.10]
  wire  _T_1281; // @[StoreQueue.scala 103:75:@420.10]
  wire  _T_1282; // @[StoreQueue.scala 103:49:@421.10]
  wire  _T_1284; // @[StoreQueue.scala 103:9:@422.10]
  wire  _T_1285; // @[StoreQueue.scala 102:49:@423.10]
  wire  _GEN_176; // @[StoreQueue.scala 103:96:@424.10]
  wire  _GEN_177; // @[StoreQueue.scala 100:102:@414.8]
  wire  _GEN_178; // @[StoreQueue.scala 98:26:@407.6]
  wire  _GEN_179; // @[StoreQueue.scala 94:35:@392.4]
  wire [3:0] _T_1298; // @[util.scala 10:8:@435.6]
  wire [3:0] _GEN_27; // @[util.scala 10:14:@436.6]
  wire [3:0] _T_1299; // @[util.scala 10:14:@436.6]
  wire  _T_1300; // @[StoreQueue.scala 96:56:@437.6]
  wire  _T_1301; // @[StoreQueue.scala 95:50:@438.6]
  wire  _T_1303; // @[StoreQueue.scala 95:35:@439.6]
  wire  _T_1305; // @[StoreQueue.scala 100:35:@447.8]
  wire  _T_1306; // @[StoreQueue.scala 100:87:@448.8]
  wire  _T_1307; // @[StoreQueue.scala 100:61:@449.8]
  wire  _T_1310; // @[StoreQueue.scala 103:23:@455.10]
  wire  _T_1311; // @[StoreQueue.scala 103:75:@456.10]
  wire  _T_1312; // @[StoreQueue.scala 103:49:@457.10]
  wire  _T_1314; // @[StoreQueue.scala 103:9:@458.10]
  wire  _T_1315; // @[StoreQueue.scala 102:49:@459.10]
  wire  _GEN_188; // @[StoreQueue.scala 103:96:@460.10]
  wire  _GEN_189; // @[StoreQueue.scala 100:102:@450.8]
  wire  _GEN_190; // @[StoreQueue.scala 98:26:@443.6]
  wire  _GEN_191; // @[StoreQueue.scala 94:35:@428.4]
  wire [3:0] _T_1328; // @[util.scala 10:8:@471.6]
  wire [3:0] _GEN_28; // @[util.scala 10:14:@472.6]
  wire [3:0] _T_1329; // @[util.scala 10:14:@472.6]
  wire  _T_1330; // @[StoreQueue.scala 96:56:@473.6]
  wire  _T_1331; // @[StoreQueue.scala 95:50:@474.6]
  wire  _T_1333; // @[StoreQueue.scala 95:35:@475.6]
  wire  _T_1335; // @[StoreQueue.scala 100:35:@483.8]
  wire  _T_1336; // @[StoreQueue.scala 100:87:@484.8]
  wire  _T_1337; // @[StoreQueue.scala 100:61:@485.8]
  wire  _T_1340; // @[StoreQueue.scala 103:23:@491.10]
  wire  _T_1341; // @[StoreQueue.scala 103:75:@492.10]
  wire  _T_1342; // @[StoreQueue.scala 103:49:@493.10]
  wire  _T_1344; // @[StoreQueue.scala 103:9:@494.10]
  wire  _T_1345; // @[StoreQueue.scala 102:49:@495.10]
  wire  _GEN_200; // @[StoreQueue.scala 103:96:@496.10]
  wire  _GEN_201; // @[StoreQueue.scala 100:102:@486.8]
  wire  _GEN_202; // @[StoreQueue.scala 98:26:@479.6]
  wire  _GEN_203; // @[StoreQueue.scala 94:35:@464.4]
  wire [3:0] _T_1358; // @[util.scala 10:8:@507.6]
  wire [3:0] _GEN_29; // @[util.scala 10:14:@508.6]
  wire [3:0] _T_1359; // @[util.scala 10:14:@508.6]
  wire  _T_1360; // @[StoreQueue.scala 96:56:@509.6]
  wire  _T_1361; // @[StoreQueue.scala 95:50:@510.6]
  wire  _T_1363; // @[StoreQueue.scala 95:35:@511.6]
  wire  _T_1365; // @[StoreQueue.scala 100:35:@519.8]
  wire  _T_1366; // @[StoreQueue.scala 100:87:@520.8]
  wire  _T_1367; // @[StoreQueue.scala 100:61:@521.8]
  wire  _T_1370; // @[StoreQueue.scala 103:23:@527.10]
  wire  _T_1371; // @[StoreQueue.scala 103:75:@528.10]
  wire  _T_1372; // @[StoreQueue.scala 103:49:@529.10]
  wire  _T_1374; // @[StoreQueue.scala 103:9:@530.10]
  wire  _T_1375; // @[StoreQueue.scala 102:49:@531.10]
  wire  _GEN_212; // @[StoreQueue.scala 103:96:@532.10]
  wire  _GEN_213; // @[StoreQueue.scala 100:102:@522.8]
  wire  _GEN_214; // @[StoreQueue.scala 98:26:@515.6]
  wire  _GEN_215; // @[StoreQueue.scala 94:35:@500.4]
  wire [3:0] _T_1388; // @[util.scala 10:8:@543.6]
  wire [3:0] _GEN_30; // @[util.scala 10:14:@544.6]
  wire [3:0] _T_1389; // @[util.scala 10:14:@544.6]
  wire  _T_1390; // @[StoreQueue.scala 96:56:@545.6]
  wire  _T_1391; // @[StoreQueue.scala 95:50:@546.6]
  wire  _T_1393; // @[StoreQueue.scala 95:35:@547.6]
  wire  _T_1395; // @[StoreQueue.scala 100:35:@555.8]
  wire  _T_1396; // @[StoreQueue.scala 100:87:@556.8]
  wire  _T_1397; // @[StoreQueue.scala 100:61:@557.8]
  wire  _T_1400; // @[StoreQueue.scala 103:23:@563.10]
  wire  _T_1401; // @[StoreQueue.scala 103:75:@564.10]
  wire  _T_1402; // @[StoreQueue.scala 103:49:@565.10]
  wire  _T_1404; // @[StoreQueue.scala 103:9:@566.10]
  wire  _T_1405; // @[StoreQueue.scala 102:49:@567.10]
  wire  _GEN_224; // @[StoreQueue.scala 103:96:@568.10]
  wire  _GEN_225; // @[StoreQueue.scala 100:102:@558.8]
  wire  _GEN_226; // @[StoreQueue.scala 98:26:@551.6]
  wire  _GEN_227; // @[StoreQueue.scala 94:35:@536.4]
  wire [3:0] _T_1418; // @[util.scala 10:8:@579.6]
  wire [3:0] _GEN_31; // @[util.scala 10:14:@580.6]
  wire [3:0] _T_1419; // @[util.scala 10:14:@580.6]
  wire  _T_1420; // @[StoreQueue.scala 96:56:@581.6]
  wire  _T_1421; // @[StoreQueue.scala 95:50:@582.6]
  wire  _T_1423; // @[StoreQueue.scala 95:35:@583.6]
  wire  _T_1425; // @[StoreQueue.scala 100:35:@591.8]
  wire  _T_1426; // @[StoreQueue.scala 100:87:@592.8]
  wire  _T_1427; // @[StoreQueue.scala 100:61:@593.8]
  wire  _T_1430; // @[StoreQueue.scala 103:23:@599.10]
  wire  _T_1431; // @[StoreQueue.scala 103:75:@600.10]
  wire  _T_1432; // @[StoreQueue.scala 103:49:@601.10]
  wire  _T_1434; // @[StoreQueue.scala 103:9:@602.10]
  wire  _T_1435; // @[StoreQueue.scala 102:49:@603.10]
  wire  _GEN_236; // @[StoreQueue.scala 103:96:@604.10]
  wire  _GEN_237; // @[StoreQueue.scala 100:102:@594.8]
  wire  _GEN_238; // @[StoreQueue.scala 98:26:@587.6]
  wire  _GEN_239; // @[StoreQueue.scala 94:35:@572.4]
  wire  _T_1437; // @[StoreQueue.scala 119:103:@608.4]
  wire  _T_1439; // @[StoreQueue.scala 120:17:@609.4]
  wire  _T_1441; // @[StoreQueue.scala 120:35:@610.4]
  wire  _T_1442; // @[StoreQueue.scala 120:26:@611.4]
  wire  _T_1444; // @[StoreQueue.scala 120:50:@612.4]
  wire  _T_1446; // @[StoreQueue.scala 120:81:@613.4]
  wire  _T_1448; // @[StoreQueue.scala 120:99:@614.4]
  wire  _T_1449; // @[StoreQueue.scala 120:90:@615.4]
  wire  _T_1451; // @[StoreQueue.scala 120:67:@616.4]
  wire  _T_1452; // @[StoreQueue.scala 120:64:@617.4]
  wire  validEntriesInLoadQ_0; // @[StoreQueue.scala 119:90:@618.4]
  wire  _T_1456; // @[StoreQueue.scala 120:17:@620.4]
  wire  _T_1458; // @[StoreQueue.scala 120:35:@621.4]
  wire  _T_1459; // @[StoreQueue.scala 120:26:@622.4]
  wire  _T_1463; // @[StoreQueue.scala 120:81:@624.4]
  wire  _T_1465; // @[StoreQueue.scala 120:99:@625.4]
  wire  _T_1466; // @[StoreQueue.scala 120:90:@626.4]
  wire  _T_1468; // @[StoreQueue.scala 120:67:@627.4]
  wire  _T_1469; // @[StoreQueue.scala 120:64:@628.4]
  wire  validEntriesInLoadQ_1; // @[StoreQueue.scala 119:90:@629.4]
  wire  _T_1473; // @[StoreQueue.scala 120:17:@631.4]
  wire  _T_1475; // @[StoreQueue.scala 120:35:@632.4]
  wire  _T_1476; // @[StoreQueue.scala 120:26:@633.4]
  wire  _T_1480; // @[StoreQueue.scala 120:81:@635.4]
  wire  _T_1482; // @[StoreQueue.scala 120:99:@636.4]
  wire  _T_1483; // @[StoreQueue.scala 120:90:@637.4]
  wire  _T_1485; // @[StoreQueue.scala 120:67:@638.4]
  wire  _T_1486; // @[StoreQueue.scala 120:64:@639.4]
  wire  validEntriesInLoadQ_2; // @[StoreQueue.scala 119:90:@640.4]
  wire  _T_1490; // @[StoreQueue.scala 120:17:@642.4]
  wire  _T_1492; // @[StoreQueue.scala 120:35:@643.4]
  wire  _T_1493; // @[StoreQueue.scala 120:26:@644.4]
  wire  _T_1497; // @[StoreQueue.scala 120:81:@646.4]
  wire  _T_1499; // @[StoreQueue.scala 120:99:@647.4]
  wire  _T_1500; // @[StoreQueue.scala 120:90:@648.4]
  wire  _T_1502; // @[StoreQueue.scala 120:67:@649.4]
  wire  _T_1503; // @[StoreQueue.scala 120:64:@650.4]
  wire  validEntriesInLoadQ_3; // @[StoreQueue.scala 119:90:@651.4]
  wire  _T_1507; // @[StoreQueue.scala 120:17:@653.4]
  wire  _T_1509; // @[StoreQueue.scala 120:35:@654.4]
  wire  _T_1510; // @[StoreQueue.scala 120:26:@655.4]
  wire  _T_1514; // @[StoreQueue.scala 120:81:@657.4]
  wire  _T_1516; // @[StoreQueue.scala 120:99:@658.4]
  wire  _T_1517; // @[StoreQueue.scala 120:90:@659.4]
  wire  _T_1519; // @[StoreQueue.scala 120:67:@660.4]
  wire  _T_1520; // @[StoreQueue.scala 120:64:@661.4]
  wire  validEntriesInLoadQ_4; // @[StoreQueue.scala 119:90:@662.4]
  wire  _T_1524; // @[StoreQueue.scala 120:17:@664.4]
  wire  _T_1526; // @[StoreQueue.scala 120:35:@665.4]
  wire  _T_1527; // @[StoreQueue.scala 120:26:@666.4]
  wire  _T_1531; // @[StoreQueue.scala 120:81:@668.4]
  wire  _T_1533; // @[StoreQueue.scala 120:99:@669.4]
  wire  _T_1534; // @[StoreQueue.scala 120:90:@670.4]
  wire  _T_1536; // @[StoreQueue.scala 120:67:@671.4]
  wire  _T_1537; // @[StoreQueue.scala 120:64:@672.4]
  wire  validEntriesInLoadQ_5; // @[StoreQueue.scala 119:90:@673.4]
  wire  _T_1541; // @[StoreQueue.scala 120:17:@675.4]
  wire  _T_1543; // @[StoreQueue.scala 120:35:@676.4]
  wire  _T_1544; // @[StoreQueue.scala 120:26:@677.4]
  wire  _T_1548; // @[StoreQueue.scala 120:81:@679.4]
  wire  _T_1550; // @[StoreQueue.scala 120:99:@680.4]
  wire  _T_1551; // @[StoreQueue.scala 120:90:@681.4]
  wire  _T_1553; // @[StoreQueue.scala 120:67:@682.4]
  wire  _T_1554; // @[StoreQueue.scala 120:64:@683.4]
  wire  validEntriesInLoadQ_6; // @[StoreQueue.scala 119:90:@684.4]
  wire  validEntriesInLoadQ_7; // @[StoreQueue.scala 119:90:@695.4]
  wire [2:0] _GEN_241; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_242; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_243; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_244; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_245; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_246; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_247; // @[StoreQueue.scala 126:96:@705.4]
  wire  _T_1589; // @[StoreQueue.scala 126:96:@705.4]
  wire  loadsToCheck_0; // @[StoreQueue.scala 126:83:@713.4]
  wire  _T_1619; // @[StoreQueue.scala 127:37:@716.4]
  wire  _T_1620; // @[StoreQueue.scala 127:28:@717.4]
  wire  _T_1625; // @[StoreQueue.scala 127:71:@718.4]
  wire  _T_1628; // @[StoreQueue.scala 127:79:@720.4]
  wire  _T_1630; // @[StoreQueue.scala 127:55:@721.4]
  wire  loadsToCheck_1; // @[StoreQueue.scala 126:83:@722.4]
  wire  _T_1642; // @[StoreQueue.scala 127:37:@725.4]
  wire  _T_1643; // @[StoreQueue.scala 127:28:@726.4]
  wire  _T_1648; // @[StoreQueue.scala 127:71:@727.4]
  wire  _T_1651; // @[StoreQueue.scala 127:79:@729.4]
  wire  _T_1653; // @[StoreQueue.scala 127:55:@730.4]
  wire  loadsToCheck_2; // @[StoreQueue.scala 126:83:@731.4]
  wire  _T_1665; // @[StoreQueue.scala 127:37:@734.4]
  wire  _T_1666; // @[StoreQueue.scala 127:28:@735.4]
  wire  _T_1671; // @[StoreQueue.scala 127:71:@736.4]
  wire  _T_1674; // @[StoreQueue.scala 127:79:@738.4]
  wire  _T_1676; // @[StoreQueue.scala 127:55:@739.4]
  wire  loadsToCheck_3; // @[StoreQueue.scala 126:83:@740.4]
  wire  _T_1688; // @[StoreQueue.scala 127:37:@743.4]
  wire  _T_1689; // @[StoreQueue.scala 127:28:@744.4]
  wire  _T_1694; // @[StoreQueue.scala 127:71:@745.4]
  wire  _T_1697; // @[StoreQueue.scala 127:79:@747.4]
  wire  _T_1699; // @[StoreQueue.scala 127:55:@748.4]
  wire  loadsToCheck_4; // @[StoreQueue.scala 126:83:@749.4]
  wire  _T_1711; // @[StoreQueue.scala 127:37:@752.4]
  wire  _T_1712; // @[StoreQueue.scala 127:28:@753.4]
  wire  _T_1717; // @[StoreQueue.scala 127:71:@754.4]
  wire  _T_1720; // @[StoreQueue.scala 127:79:@756.4]
  wire  _T_1722; // @[StoreQueue.scala 127:55:@757.4]
  wire  loadsToCheck_5; // @[StoreQueue.scala 126:83:@758.4]
  wire  _T_1734; // @[StoreQueue.scala 127:37:@761.4]
  wire  _T_1735; // @[StoreQueue.scala 127:28:@762.4]
  wire  _T_1740; // @[StoreQueue.scala 127:71:@763.4]
  wire  _T_1743; // @[StoreQueue.scala 127:79:@765.4]
  wire  _T_1745; // @[StoreQueue.scala 127:55:@766.4]
  wire  loadsToCheck_6; // @[StoreQueue.scala 126:83:@767.4]
  wire  _T_1757; // @[StoreQueue.scala 127:37:@770.4]
  wire  loadsToCheck_7; // @[StoreQueue.scala 126:83:@776.4]
  wire  _T_1783; // @[StoreQueue.scala 133:16:@786.4]
  wire  _GEN_249; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_250; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_251; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_252; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_253; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_254; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_255; // @[StoreQueue.scala 133:24:@787.4]
  wire  entriesToCheck_0; // @[StoreQueue.scala 133:24:@787.4]
  wire  _T_1788; // @[StoreQueue.scala 133:16:@788.4]
  wire  entriesToCheck_1; // @[StoreQueue.scala 133:24:@789.4]
  wire  _T_1793; // @[StoreQueue.scala 133:16:@790.4]
  wire  entriesToCheck_2; // @[StoreQueue.scala 133:24:@791.4]
  wire  _T_1798; // @[StoreQueue.scala 133:16:@792.4]
  wire  entriesToCheck_3; // @[StoreQueue.scala 133:24:@793.4]
  wire  _T_1803; // @[StoreQueue.scala 133:16:@794.4]
  wire  entriesToCheck_4; // @[StoreQueue.scala 133:24:@795.4]
  wire  _T_1808; // @[StoreQueue.scala 133:16:@796.4]
  wire  entriesToCheck_5; // @[StoreQueue.scala 133:24:@797.4]
  wire  _T_1813; // @[StoreQueue.scala 133:16:@798.4]
  wire  entriesToCheck_6; // @[StoreQueue.scala 133:24:@799.4]
  wire  _T_1818; // @[StoreQueue.scala 133:16:@800.4]
  wire  entriesToCheck_7; // @[StoreQueue.scala 133:24:@801.4]
  wire  _T_1850; // @[StoreQueue.scala 140:34:@812.4]
  wire  _T_1851; // @[StoreQueue.scala 140:64:@813.4]
  wire [31:0] _GEN_257; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_258; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_259; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_260; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_261; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_262; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_263; // @[StoreQueue.scala 141:51:@814.4]
  wire  _T_1855; // @[StoreQueue.scala 141:51:@814.4]
  wire  _T_1856; // @[StoreQueue.scala 141:36:@815.4]
  wire  noConflicts_0; // @[StoreQueue.scala 140:95:@816.4]
  wire  _T_1859; // @[StoreQueue.scala 140:34:@818.4]
  wire  _T_1860; // @[StoreQueue.scala 140:64:@819.4]
  wire  _T_1864; // @[StoreQueue.scala 141:51:@820.4]
  wire  _T_1865; // @[StoreQueue.scala 141:36:@821.4]
  wire  noConflicts_1; // @[StoreQueue.scala 140:95:@822.4]
  wire  _T_1868; // @[StoreQueue.scala 140:34:@824.4]
  wire  _T_1869; // @[StoreQueue.scala 140:64:@825.4]
  wire  _T_1873; // @[StoreQueue.scala 141:51:@826.4]
  wire  _T_1874; // @[StoreQueue.scala 141:36:@827.4]
  wire  noConflicts_2; // @[StoreQueue.scala 140:95:@828.4]
  wire  _T_1877; // @[StoreQueue.scala 140:34:@830.4]
  wire  _T_1878; // @[StoreQueue.scala 140:64:@831.4]
  wire  _T_1882; // @[StoreQueue.scala 141:51:@832.4]
  wire  _T_1883; // @[StoreQueue.scala 141:36:@833.4]
  wire  noConflicts_3; // @[StoreQueue.scala 140:95:@834.4]
  wire  _T_1886; // @[StoreQueue.scala 140:34:@836.4]
  wire  _T_1887; // @[StoreQueue.scala 140:64:@837.4]
  wire  _T_1891; // @[StoreQueue.scala 141:51:@838.4]
  wire  _T_1892; // @[StoreQueue.scala 141:36:@839.4]
  wire  noConflicts_4; // @[StoreQueue.scala 140:95:@840.4]
  wire  _T_1895; // @[StoreQueue.scala 140:34:@842.4]
  wire  _T_1896; // @[StoreQueue.scala 140:64:@843.4]
  wire  _T_1900; // @[StoreQueue.scala 141:51:@844.4]
  wire  _T_1901; // @[StoreQueue.scala 141:36:@845.4]
  wire  noConflicts_5; // @[StoreQueue.scala 140:95:@846.4]
  wire  _T_1904; // @[StoreQueue.scala 140:34:@848.4]
  wire  _T_1905; // @[StoreQueue.scala 140:64:@849.4]
  wire  _T_1909; // @[StoreQueue.scala 141:51:@850.4]
  wire  _T_1910; // @[StoreQueue.scala 141:36:@851.4]
  wire  noConflicts_6; // @[StoreQueue.scala 140:95:@852.4]
  wire  _T_1913; // @[StoreQueue.scala 140:34:@854.4]
  wire  _T_1914; // @[StoreQueue.scala 140:64:@855.4]
  wire  _T_1918; // @[StoreQueue.scala 141:51:@856.4]
  wire  _T_1919; // @[StoreQueue.scala 141:36:@857.4]
  wire  noConflicts_7; // @[StoreQueue.scala 140:95:@858.4]
  wire  _GEN_265; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_266; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_267; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_268; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_269; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_270; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_271; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_273; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_274; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_275; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_276; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_277; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_278; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_279; // @[StoreQueue.scala 154:44:@860.4]
  wire  _T_1927; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_281; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_282; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_283; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_284; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_285; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_286; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_287; // @[StoreQueue.scala 154:66:@861.4]
  wire  _T_1932; // @[StoreQueue.scala 154:66:@861.4]
  wire  _T_1933; // @[StoreQueue.scala 154:63:@862.4]
  wire  _T_1936; // @[StoreQueue.scala 154:109:@864.4]
  wire  _T_1937; // @[StoreQueue.scala 154:109:@865.4]
  wire  _T_1938; // @[StoreQueue.scala 154:109:@866.4]
  wire  _T_1939; // @[StoreQueue.scala 154:109:@867.4]
  wire  _T_1940; // @[StoreQueue.scala 154:109:@868.4]
  wire  _T_1941; // @[StoreQueue.scala 154:109:@869.4]
  wire  _T_1942; // @[StoreQueue.scala 154:109:@870.4]
  wire  storeRequest; // @[StoreQueue.scala 154:88:@871.4]
  wire  _T_1945; // @[StoreQueue.scala 164:23:@876.6]
  wire  _T_1946; // @[StoreQueue.scala 164:43:@877.6]
  wire  _T_1947; // @[StoreQueue.scala 164:59:@878.6]
  wire  _GEN_288; // @[StoreQueue.scala 164:86:@879.6]
  wire  _GEN_289; // @[StoreQueue.scala 162:37:@872.4]
  wire  _T_1951; // @[StoreQueue.scala 164:23:@886.6]
  wire  _T_1952; // @[StoreQueue.scala 164:43:@887.6]
  wire  _T_1953; // @[StoreQueue.scala 164:59:@888.6]
  wire  _GEN_290; // @[StoreQueue.scala 164:86:@889.6]
  wire  _GEN_291; // @[StoreQueue.scala 162:37:@882.4]
  wire  _T_1957; // @[StoreQueue.scala 164:23:@896.6]
  wire  _T_1958; // @[StoreQueue.scala 164:43:@897.6]
  wire  _T_1959; // @[StoreQueue.scala 164:59:@898.6]
  wire  _GEN_292; // @[StoreQueue.scala 164:86:@899.6]
  wire  _GEN_293; // @[StoreQueue.scala 162:37:@892.4]
  wire  _T_1963; // @[StoreQueue.scala 164:23:@906.6]
  wire  _T_1964; // @[StoreQueue.scala 164:43:@907.6]
  wire  _T_1965; // @[StoreQueue.scala 164:59:@908.6]
  wire  _GEN_294; // @[StoreQueue.scala 164:86:@909.6]
  wire  _GEN_295; // @[StoreQueue.scala 162:37:@902.4]
  wire  _T_1969; // @[StoreQueue.scala 164:23:@916.6]
  wire  _T_1970; // @[StoreQueue.scala 164:43:@917.6]
  wire  _T_1971; // @[StoreQueue.scala 164:59:@918.6]
  wire  _GEN_296; // @[StoreQueue.scala 164:86:@919.6]
  wire  _GEN_297; // @[StoreQueue.scala 162:37:@912.4]
  wire  _T_1975; // @[StoreQueue.scala 164:23:@926.6]
  wire  _T_1976; // @[StoreQueue.scala 164:43:@927.6]
  wire  _T_1977; // @[StoreQueue.scala 164:59:@928.6]
  wire  _GEN_298; // @[StoreQueue.scala 164:86:@929.6]
  wire  _GEN_299; // @[StoreQueue.scala 162:37:@922.4]
  wire  _T_1981; // @[StoreQueue.scala 164:23:@936.6]
  wire  _T_1982; // @[StoreQueue.scala 164:43:@937.6]
  wire  _T_1983; // @[StoreQueue.scala 164:59:@938.6]
  wire  _GEN_300; // @[StoreQueue.scala 164:86:@939.6]
  wire  _GEN_301; // @[StoreQueue.scala 162:37:@932.4]
  wire  _T_1987; // @[StoreQueue.scala 164:23:@946.6]
  wire  _T_1988; // @[StoreQueue.scala 164:43:@947.6]
  wire  _T_1989; // @[StoreQueue.scala 164:59:@948.6]
  wire  _GEN_302; // @[StoreQueue.scala 164:86:@949.6]
  wire  _GEN_303; // @[StoreQueue.scala 162:37:@942.4]
  wire  entriesPorts_0_0; // @[StoreQueue.scala 180:72:@953.4]
  wire  entriesPorts_0_1; // @[StoreQueue.scala 180:72:@955.4]
  wire  entriesPorts_0_2; // @[StoreQueue.scala 180:72:@957.4]
  wire  entriesPorts_0_3; // @[StoreQueue.scala 180:72:@959.4]
  wire  entriesPorts_0_4; // @[StoreQueue.scala 180:72:@961.4]
  wire  entriesPorts_0_5; // @[StoreQueue.scala 180:72:@963.4]
  wire  entriesPorts_0_6; // @[StoreQueue.scala 180:72:@965.4]
  wire  entriesPorts_0_7; // @[StoreQueue.scala 180:72:@967.4]
  wire  _T_2266; // @[StoreQueue.scala 192:91:@971.4]
  wire  _T_2267; // @[StoreQueue.scala 192:88:@972.4]
  wire  _T_2269; // @[StoreQueue.scala 192:91:@973.4]
  wire  _T_2270; // @[StoreQueue.scala 192:88:@974.4]
  wire  _T_2272; // @[StoreQueue.scala 192:91:@975.4]
  wire  _T_2273; // @[StoreQueue.scala 192:88:@976.4]
  wire  _T_2275; // @[StoreQueue.scala 192:91:@977.4]
  wire  _T_2276; // @[StoreQueue.scala 192:88:@978.4]
  wire  _T_2278; // @[StoreQueue.scala 192:91:@979.4]
  wire  _T_2279; // @[StoreQueue.scala 192:88:@980.4]
  wire  _T_2281; // @[StoreQueue.scala 192:91:@981.4]
  wire  _T_2282; // @[StoreQueue.scala 192:88:@982.4]
  wire  _T_2284; // @[StoreQueue.scala 192:91:@983.4]
  wire  _T_2285; // @[StoreQueue.scala 192:88:@984.4]
  wire  _T_2287; // @[StoreQueue.scala 192:91:@985.4]
  wire  _T_2288; // @[StoreQueue.scala 192:88:@986.4]
  wire  _T_2304; // @[StoreQueue.scala 193:91:@996.4]
  wire  _T_2305; // @[StoreQueue.scala 193:88:@997.4]
  wire  _T_2307; // @[StoreQueue.scala 193:91:@998.4]
  wire  _T_2308; // @[StoreQueue.scala 193:88:@999.4]
  wire  _T_2310; // @[StoreQueue.scala 193:91:@1000.4]
  wire  _T_2311; // @[StoreQueue.scala 193:88:@1001.4]
  wire  _T_2313; // @[StoreQueue.scala 193:91:@1002.4]
  wire  _T_2314; // @[StoreQueue.scala 193:88:@1003.4]
  wire  _T_2316; // @[StoreQueue.scala 193:91:@1004.4]
  wire  _T_2317; // @[StoreQueue.scala 193:88:@1005.4]
  wire  _T_2319; // @[StoreQueue.scala 193:91:@1006.4]
  wire  _T_2320; // @[StoreQueue.scala 193:88:@1007.4]
  wire  _T_2322; // @[StoreQueue.scala 193:91:@1008.4]
  wire  _T_2323; // @[StoreQueue.scala 193:88:@1009.4]
  wire  _T_2325; // @[StoreQueue.scala 193:91:@1010.4]
  wire  _T_2326; // @[StoreQueue.scala 193:88:@1011.4]
  wire [7:0] _T_2343; // @[OneHot.scala 52:12:@1022.4]
  wire  _T_2345; // @[util.scala 33:60:@1024.4]
  wire  _T_2346; // @[util.scala 33:60:@1025.4]
  wire  _T_2347; // @[util.scala 33:60:@1026.4]
  wire  _T_2348; // @[util.scala 33:60:@1027.4]
  wire  _T_2349; // @[util.scala 33:60:@1028.4]
  wire  _T_2350; // @[util.scala 33:60:@1029.4]
  wire  _T_2351; // @[util.scala 33:60:@1030.4]
  wire  _T_2352; // @[util.scala 33:60:@1031.4]
  wire [7:0] _T_2377; // @[Mux.scala 31:69:@1041.4]
  wire [7:0] _T_2378; // @[Mux.scala 31:69:@1042.4]
  wire [7:0] _T_2379; // @[Mux.scala 31:69:@1043.4]
  wire [7:0] _T_2380; // @[Mux.scala 31:69:@1044.4]
  wire [7:0] _T_2381; // @[Mux.scala 31:69:@1045.4]
  wire [7:0] _T_2382; // @[Mux.scala 31:69:@1046.4]
  wire [7:0] _T_2383; // @[Mux.scala 31:69:@1047.4]
  wire [7:0] _T_2384; // @[Mux.scala 31:69:@1048.4]
  wire  _T_2385; // @[OneHot.scala 66:30:@1049.4]
  wire  _T_2386; // @[OneHot.scala 66:30:@1050.4]
  wire  _T_2387; // @[OneHot.scala 66:30:@1051.4]
  wire  _T_2388; // @[OneHot.scala 66:30:@1052.4]
  wire  _T_2389; // @[OneHot.scala 66:30:@1053.4]
  wire  _T_2390; // @[OneHot.scala 66:30:@1054.4]
  wire  _T_2391; // @[OneHot.scala 66:30:@1055.4]
  wire  _T_2392; // @[OneHot.scala 66:30:@1056.4]
  wire [7:0] _T_2417; // @[Mux.scala 31:69:@1066.4]
  wire [7:0] _T_2418; // @[Mux.scala 31:69:@1067.4]
  wire [7:0] _T_2419; // @[Mux.scala 31:69:@1068.4]
  wire [7:0] _T_2420; // @[Mux.scala 31:69:@1069.4]
  wire [7:0] _T_2421; // @[Mux.scala 31:69:@1070.4]
  wire [7:0] _T_2422; // @[Mux.scala 31:69:@1071.4]
  wire [7:0] _T_2423; // @[Mux.scala 31:69:@1072.4]
  wire [7:0] _T_2424; // @[Mux.scala 31:69:@1073.4]
  wire  _T_2425; // @[OneHot.scala 66:30:@1074.4]
  wire  _T_2426; // @[OneHot.scala 66:30:@1075.4]
  wire  _T_2427; // @[OneHot.scala 66:30:@1076.4]
  wire  _T_2428; // @[OneHot.scala 66:30:@1077.4]
  wire  _T_2429; // @[OneHot.scala 66:30:@1078.4]
  wire  _T_2430; // @[OneHot.scala 66:30:@1079.4]
  wire  _T_2431; // @[OneHot.scala 66:30:@1080.4]
  wire  _T_2432; // @[OneHot.scala 66:30:@1081.4]
  wire [7:0] _T_2457; // @[Mux.scala 31:69:@1091.4]
  wire [7:0] _T_2458; // @[Mux.scala 31:69:@1092.4]
  wire [7:0] _T_2459; // @[Mux.scala 31:69:@1093.4]
  wire [7:0] _T_2460; // @[Mux.scala 31:69:@1094.4]
  wire [7:0] _T_2461; // @[Mux.scala 31:69:@1095.4]
  wire [7:0] _T_2462; // @[Mux.scala 31:69:@1096.4]
  wire [7:0] _T_2463; // @[Mux.scala 31:69:@1097.4]
  wire [7:0] _T_2464; // @[Mux.scala 31:69:@1098.4]
  wire  _T_2465; // @[OneHot.scala 66:30:@1099.4]
  wire  _T_2466; // @[OneHot.scala 66:30:@1100.4]
  wire  _T_2467; // @[OneHot.scala 66:30:@1101.4]
  wire  _T_2468; // @[OneHot.scala 66:30:@1102.4]
  wire  _T_2469; // @[OneHot.scala 66:30:@1103.4]
  wire  _T_2470; // @[OneHot.scala 66:30:@1104.4]
  wire  _T_2471; // @[OneHot.scala 66:30:@1105.4]
  wire  _T_2472; // @[OneHot.scala 66:30:@1106.4]
  wire [7:0] _T_2497; // @[Mux.scala 31:69:@1116.4]
  wire [7:0] _T_2498; // @[Mux.scala 31:69:@1117.4]
  wire [7:0] _T_2499; // @[Mux.scala 31:69:@1118.4]
  wire [7:0] _T_2500; // @[Mux.scala 31:69:@1119.4]
  wire [7:0] _T_2501; // @[Mux.scala 31:69:@1120.4]
  wire [7:0] _T_2502; // @[Mux.scala 31:69:@1121.4]
  wire [7:0] _T_2503; // @[Mux.scala 31:69:@1122.4]
  wire [7:0] _T_2504; // @[Mux.scala 31:69:@1123.4]
  wire  _T_2505; // @[OneHot.scala 66:30:@1124.4]
  wire  _T_2506; // @[OneHot.scala 66:30:@1125.4]
  wire  _T_2507; // @[OneHot.scala 66:30:@1126.4]
  wire  _T_2508; // @[OneHot.scala 66:30:@1127.4]
  wire  _T_2509; // @[OneHot.scala 66:30:@1128.4]
  wire  _T_2510; // @[OneHot.scala 66:30:@1129.4]
  wire  _T_2511; // @[OneHot.scala 66:30:@1130.4]
  wire  _T_2512; // @[OneHot.scala 66:30:@1131.4]
  wire [7:0] _T_2537; // @[Mux.scala 31:69:@1141.4]
  wire [7:0] _T_2538; // @[Mux.scala 31:69:@1142.4]
  wire [7:0] _T_2539; // @[Mux.scala 31:69:@1143.4]
  wire [7:0] _T_2540; // @[Mux.scala 31:69:@1144.4]
  wire [7:0] _T_2541; // @[Mux.scala 31:69:@1145.4]
  wire [7:0] _T_2542; // @[Mux.scala 31:69:@1146.4]
  wire [7:0] _T_2543; // @[Mux.scala 31:69:@1147.4]
  wire [7:0] _T_2544; // @[Mux.scala 31:69:@1148.4]
  wire  _T_2545; // @[OneHot.scala 66:30:@1149.4]
  wire  _T_2546; // @[OneHot.scala 66:30:@1150.4]
  wire  _T_2547; // @[OneHot.scala 66:30:@1151.4]
  wire  _T_2548; // @[OneHot.scala 66:30:@1152.4]
  wire  _T_2549; // @[OneHot.scala 66:30:@1153.4]
  wire  _T_2550; // @[OneHot.scala 66:30:@1154.4]
  wire  _T_2551; // @[OneHot.scala 66:30:@1155.4]
  wire  _T_2552; // @[OneHot.scala 66:30:@1156.4]
  wire [7:0] _T_2577; // @[Mux.scala 31:69:@1166.4]
  wire [7:0] _T_2578; // @[Mux.scala 31:69:@1167.4]
  wire [7:0] _T_2579; // @[Mux.scala 31:69:@1168.4]
  wire [7:0] _T_2580; // @[Mux.scala 31:69:@1169.4]
  wire [7:0] _T_2581; // @[Mux.scala 31:69:@1170.4]
  wire [7:0] _T_2582; // @[Mux.scala 31:69:@1171.4]
  wire [7:0] _T_2583; // @[Mux.scala 31:69:@1172.4]
  wire [7:0] _T_2584; // @[Mux.scala 31:69:@1173.4]
  wire  _T_2585; // @[OneHot.scala 66:30:@1174.4]
  wire  _T_2586; // @[OneHot.scala 66:30:@1175.4]
  wire  _T_2587; // @[OneHot.scala 66:30:@1176.4]
  wire  _T_2588; // @[OneHot.scala 66:30:@1177.4]
  wire  _T_2589; // @[OneHot.scala 66:30:@1178.4]
  wire  _T_2590; // @[OneHot.scala 66:30:@1179.4]
  wire  _T_2591; // @[OneHot.scala 66:30:@1180.4]
  wire  _T_2592; // @[OneHot.scala 66:30:@1181.4]
  wire [7:0] _T_2617; // @[Mux.scala 31:69:@1191.4]
  wire [7:0] _T_2618; // @[Mux.scala 31:69:@1192.4]
  wire [7:0] _T_2619; // @[Mux.scala 31:69:@1193.4]
  wire [7:0] _T_2620; // @[Mux.scala 31:69:@1194.4]
  wire [7:0] _T_2621; // @[Mux.scala 31:69:@1195.4]
  wire [7:0] _T_2622; // @[Mux.scala 31:69:@1196.4]
  wire [7:0] _T_2623; // @[Mux.scala 31:69:@1197.4]
  wire [7:0] _T_2624; // @[Mux.scala 31:69:@1198.4]
  wire  _T_2625; // @[OneHot.scala 66:30:@1199.4]
  wire  _T_2626; // @[OneHot.scala 66:30:@1200.4]
  wire  _T_2627; // @[OneHot.scala 66:30:@1201.4]
  wire  _T_2628; // @[OneHot.scala 66:30:@1202.4]
  wire  _T_2629; // @[OneHot.scala 66:30:@1203.4]
  wire  _T_2630; // @[OneHot.scala 66:30:@1204.4]
  wire  _T_2631; // @[OneHot.scala 66:30:@1205.4]
  wire  _T_2632; // @[OneHot.scala 66:30:@1206.4]
  wire [7:0] _T_2657; // @[Mux.scala 31:69:@1216.4]
  wire [7:0] _T_2658; // @[Mux.scala 31:69:@1217.4]
  wire [7:0] _T_2659; // @[Mux.scala 31:69:@1218.4]
  wire [7:0] _T_2660; // @[Mux.scala 31:69:@1219.4]
  wire [7:0] _T_2661; // @[Mux.scala 31:69:@1220.4]
  wire [7:0] _T_2662; // @[Mux.scala 31:69:@1221.4]
  wire [7:0] _T_2663; // @[Mux.scala 31:69:@1222.4]
  wire [7:0] _T_2664; // @[Mux.scala 31:69:@1223.4]
  wire  _T_2665; // @[OneHot.scala 66:30:@1224.4]
  wire  _T_2666; // @[OneHot.scala 66:30:@1225.4]
  wire  _T_2667; // @[OneHot.scala 66:30:@1226.4]
  wire  _T_2668; // @[OneHot.scala 66:30:@1227.4]
  wire  _T_2669; // @[OneHot.scala 66:30:@1228.4]
  wire  _T_2670; // @[OneHot.scala 66:30:@1229.4]
  wire  _T_2671; // @[OneHot.scala 66:30:@1230.4]
  wire  _T_2672; // @[OneHot.scala 66:30:@1231.4]
  wire [7:0] _T_2713; // @[Mux.scala 19:72:@1247.4]
  wire [7:0] _T_2715; // @[Mux.scala 19:72:@1248.4]
  wire [7:0] _T_2722; // @[Mux.scala 19:72:@1255.4]
  wire [7:0] _T_2724; // @[Mux.scala 19:72:@1256.4]
  wire [7:0] _T_2731; // @[Mux.scala 19:72:@1263.4]
  wire [7:0] _T_2733; // @[Mux.scala 19:72:@1264.4]
  wire [7:0] _T_2740; // @[Mux.scala 19:72:@1271.4]
  wire [7:0] _T_2742; // @[Mux.scala 19:72:@1272.4]
  wire [7:0] _T_2749; // @[Mux.scala 19:72:@1279.4]
  wire [7:0] _T_2751; // @[Mux.scala 19:72:@1280.4]
  wire [7:0] _T_2758; // @[Mux.scala 19:72:@1287.4]
  wire [7:0] _T_2760; // @[Mux.scala 19:72:@1288.4]
  wire [7:0] _T_2767; // @[Mux.scala 19:72:@1295.4]
  wire [7:0] _T_2769; // @[Mux.scala 19:72:@1296.4]
  wire [7:0] _T_2776; // @[Mux.scala 19:72:@1303.4]
  wire [7:0] _T_2778; // @[Mux.scala 19:72:@1304.4]
  wire [7:0] _T_2779; // @[Mux.scala 19:72:@1305.4]
  wire [7:0] _T_2780; // @[Mux.scala 19:72:@1306.4]
  wire [7:0] _T_2781; // @[Mux.scala 19:72:@1307.4]
  wire [7:0] _T_2782; // @[Mux.scala 19:72:@1308.4]
  wire [7:0] _T_2783; // @[Mux.scala 19:72:@1309.4]
  wire [7:0] _T_2784; // @[Mux.scala 19:72:@1310.4]
  wire [7:0] _T_2785; // @[Mux.scala 19:72:@1311.4]
  wire  inputAddrPriorityPorts_0_0; // @[Mux.scala 19:72:@1315.4]
  wire  inputAddrPriorityPorts_0_1; // @[Mux.scala 19:72:@1317.4]
  wire  inputAddrPriorityPorts_0_2; // @[Mux.scala 19:72:@1319.4]
  wire  inputAddrPriorityPorts_0_3; // @[Mux.scala 19:72:@1321.4]
  wire  inputAddrPriorityPorts_0_4; // @[Mux.scala 19:72:@1323.4]
  wire  inputAddrPriorityPorts_0_5; // @[Mux.scala 19:72:@1325.4]
  wire  inputAddrPriorityPorts_0_6; // @[Mux.scala 19:72:@1327.4]
  wire  inputAddrPriorityPorts_0_7; // @[Mux.scala 19:72:@1329.4]
  wire [7:0] _T_2899; // @[Mux.scala 31:69:@1359.4]
  wire [7:0] _T_2900; // @[Mux.scala 31:69:@1360.4]
  wire [7:0] _T_2901; // @[Mux.scala 31:69:@1361.4]
  wire [7:0] _T_2902; // @[Mux.scala 31:69:@1362.4]
  wire [7:0] _T_2903; // @[Mux.scala 31:69:@1363.4]
  wire [7:0] _T_2904; // @[Mux.scala 31:69:@1364.4]
  wire [7:0] _T_2905; // @[Mux.scala 31:69:@1365.4]
  wire [7:0] _T_2906; // @[Mux.scala 31:69:@1366.4]
  wire  _T_2907; // @[OneHot.scala 66:30:@1367.4]
  wire  _T_2908; // @[OneHot.scala 66:30:@1368.4]
  wire  _T_2909; // @[OneHot.scala 66:30:@1369.4]
  wire  _T_2910; // @[OneHot.scala 66:30:@1370.4]
  wire  _T_2911; // @[OneHot.scala 66:30:@1371.4]
  wire  _T_2912; // @[OneHot.scala 66:30:@1372.4]
  wire  _T_2913; // @[OneHot.scala 66:30:@1373.4]
  wire  _T_2914; // @[OneHot.scala 66:30:@1374.4]
  wire [7:0] _T_2939; // @[Mux.scala 31:69:@1384.4]
  wire [7:0] _T_2940; // @[Mux.scala 31:69:@1385.4]
  wire [7:0] _T_2941; // @[Mux.scala 31:69:@1386.4]
  wire [7:0] _T_2942; // @[Mux.scala 31:69:@1387.4]
  wire [7:0] _T_2943; // @[Mux.scala 31:69:@1388.4]
  wire [7:0] _T_2944; // @[Mux.scala 31:69:@1389.4]
  wire [7:0] _T_2945; // @[Mux.scala 31:69:@1390.4]
  wire [7:0] _T_2946; // @[Mux.scala 31:69:@1391.4]
  wire  _T_2947; // @[OneHot.scala 66:30:@1392.4]
  wire  _T_2948; // @[OneHot.scala 66:30:@1393.4]
  wire  _T_2949; // @[OneHot.scala 66:30:@1394.4]
  wire  _T_2950; // @[OneHot.scala 66:30:@1395.4]
  wire  _T_2951; // @[OneHot.scala 66:30:@1396.4]
  wire  _T_2952; // @[OneHot.scala 66:30:@1397.4]
  wire  _T_2953; // @[OneHot.scala 66:30:@1398.4]
  wire  _T_2954; // @[OneHot.scala 66:30:@1399.4]
  wire [7:0] _T_2979; // @[Mux.scala 31:69:@1409.4]
  wire [7:0] _T_2980; // @[Mux.scala 31:69:@1410.4]
  wire [7:0] _T_2981; // @[Mux.scala 31:69:@1411.4]
  wire [7:0] _T_2982; // @[Mux.scala 31:69:@1412.4]
  wire [7:0] _T_2983; // @[Mux.scala 31:69:@1413.4]
  wire [7:0] _T_2984; // @[Mux.scala 31:69:@1414.4]
  wire [7:0] _T_2985; // @[Mux.scala 31:69:@1415.4]
  wire [7:0] _T_2986; // @[Mux.scala 31:69:@1416.4]
  wire  _T_2987; // @[OneHot.scala 66:30:@1417.4]
  wire  _T_2988; // @[OneHot.scala 66:30:@1418.4]
  wire  _T_2989; // @[OneHot.scala 66:30:@1419.4]
  wire  _T_2990; // @[OneHot.scala 66:30:@1420.4]
  wire  _T_2991; // @[OneHot.scala 66:30:@1421.4]
  wire  _T_2992; // @[OneHot.scala 66:30:@1422.4]
  wire  _T_2993; // @[OneHot.scala 66:30:@1423.4]
  wire  _T_2994; // @[OneHot.scala 66:30:@1424.4]
  wire [7:0] _T_3019; // @[Mux.scala 31:69:@1434.4]
  wire [7:0] _T_3020; // @[Mux.scala 31:69:@1435.4]
  wire [7:0] _T_3021; // @[Mux.scala 31:69:@1436.4]
  wire [7:0] _T_3022; // @[Mux.scala 31:69:@1437.4]
  wire [7:0] _T_3023; // @[Mux.scala 31:69:@1438.4]
  wire [7:0] _T_3024; // @[Mux.scala 31:69:@1439.4]
  wire [7:0] _T_3025; // @[Mux.scala 31:69:@1440.4]
  wire [7:0] _T_3026; // @[Mux.scala 31:69:@1441.4]
  wire  _T_3027; // @[OneHot.scala 66:30:@1442.4]
  wire  _T_3028; // @[OneHot.scala 66:30:@1443.4]
  wire  _T_3029; // @[OneHot.scala 66:30:@1444.4]
  wire  _T_3030; // @[OneHot.scala 66:30:@1445.4]
  wire  _T_3031; // @[OneHot.scala 66:30:@1446.4]
  wire  _T_3032; // @[OneHot.scala 66:30:@1447.4]
  wire  _T_3033; // @[OneHot.scala 66:30:@1448.4]
  wire  _T_3034; // @[OneHot.scala 66:30:@1449.4]
  wire [7:0] _T_3059; // @[Mux.scala 31:69:@1459.4]
  wire [7:0] _T_3060; // @[Mux.scala 31:69:@1460.4]
  wire [7:0] _T_3061; // @[Mux.scala 31:69:@1461.4]
  wire [7:0] _T_3062; // @[Mux.scala 31:69:@1462.4]
  wire [7:0] _T_3063; // @[Mux.scala 31:69:@1463.4]
  wire [7:0] _T_3064; // @[Mux.scala 31:69:@1464.4]
  wire [7:0] _T_3065; // @[Mux.scala 31:69:@1465.4]
  wire [7:0] _T_3066; // @[Mux.scala 31:69:@1466.4]
  wire  _T_3067; // @[OneHot.scala 66:30:@1467.4]
  wire  _T_3068; // @[OneHot.scala 66:30:@1468.4]
  wire  _T_3069; // @[OneHot.scala 66:30:@1469.4]
  wire  _T_3070; // @[OneHot.scala 66:30:@1470.4]
  wire  _T_3071; // @[OneHot.scala 66:30:@1471.4]
  wire  _T_3072; // @[OneHot.scala 66:30:@1472.4]
  wire  _T_3073; // @[OneHot.scala 66:30:@1473.4]
  wire  _T_3074; // @[OneHot.scala 66:30:@1474.4]
  wire [7:0] _T_3099; // @[Mux.scala 31:69:@1484.4]
  wire [7:0] _T_3100; // @[Mux.scala 31:69:@1485.4]
  wire [7:0] _T_3101; // @[Mux.scala 31:69:@1486.4]
  wire [7:0] _T_3102; // @[Mux.scala 31:69:@1487.4]
  wire [7:0] _T_3103; // @[Mux.scala 31:69:@1488.4]
  wire [7:0] _T_3104; // @[Mux.scala 31:69:@1489.4]
  wire [7:0] _T_3105; // @[Mux.scala 31:69:@1490.4]
  wire [7:0] _T_3106; // @[Mux.scala 31:69:@1491.4]
  wire  _T_3107; // @[OneHot.scala 66:30:@1492.4]
  wire  _T_3108; // @[OneHot.scala 66:30:@1493.4]
  wire  _T_3109; // @[OneHot.scala 66:30:@1494.4]
  wire  _T_3110; // @[OneHot.scala 66:30:@1495.4]
  wire  _T_3111; // @[OneHot.scala 66:30:@1496.4]
  wire  _T_3112; // @[OneHot.scala 66:30:@1497.4]
  wire  _T_3113; // @[OneHot.scala 66:30:@1498.4]
  wire  _T_3114; // @[OneHot.scala 66:30:@1499.4]
  wire [7:0] _T_3139; // @[Mux.scala 31:69:@1509.4]
  wire [7:0] _T_3140; // @[Mux.scala 31:69:@1510.4]
  wire [7:0] _T_3141; // @[Mux.scala 31:69:@1511.4]
  wire [7:0] _T_3142; // @[Mux.scala 31:69:@1512.4]
  wire [7:0] _T_3143; // @[Mux.scala 31:69:@1513.4]
  wire [7:0] _T_3144; // @[Mux.scala 31:69:@1514.4]
  wire [7:0] _T_3145; // @[Mux.scala 31:69:@1515.4]
  wire [7:0] _T_3146; // @[Mux.scala 31:69:@1516.4]
  wire  _T_3147; // @[OneHot.scala 66:30:@1517.4]
  wire  _T_3148; // @[OneHot.scala 66:30:@1518.4]
  wire  _T_3149; // @[OneHot.scala 66:30:@1519.4]
  wire  _T_3150; // @[OneHot.scala 66:30:@1520.4]
  wire  _T_3151; // @[OneHot.scala 66:30:@1521.4]
  wire  _T_3152; // @[OneHot.scala 66:30:@1522.4]
  wire  _T_3153; // @[OneHot.scala 66:30:@1523.4]
  wire  _T_3154; // @[OneHot.scala 66:30:@1524.4]
  wire [7:0] _T_3179; // @[Mux.scala 31:69:@1534.4]
  wire [7:0] _T_3180; // @[Mux.scala 31:69:@1535.4]
  wire [7:0] _T_3181; // @[Mux.scala 31:69:@1536.4]
  wire [7:0] _T_3182; // @[Mux.scala 31:69:@1537.4]
  wire [7:0] _T_3183; // @[Mux.scala 31:69:@1538.4]
  wire [7:0] _T_3184; // @[Mux.scala 31:69:@1539.4]
  wire [7:0] _T_3185; // @[Mux.scala 31:69:@1540.4]
  wire [7:0] _T_3186; // @[Mux.scala 31:69:@1541.4]
  wire  _T_3187; // @[OneHot.scala 66:30:@1542.4]
  wire  _T_3188; // @[OneHot.scala 66:30:@1543.4]
  wire  _T_3189; // @[OneHot.scala 66:30:@1544.4]
  wire  _T_3190; // @[OneHot.scala 66:30:@1545.4]
  wire  _T_3191; // @[OneHot.scala 66:30:@1546.4]
  wire  _T_3192; // @[OneHot.scala 66:30:@1547.4]
  wire  _T_3193; // @[OneHot.scala 66:30:@1548.4]
  wire  _T_3194; // @[OneHot.scala 66:30:@1549.4]
  wire [7:0] _T_3235; // @[Mux.scala 19:72:@1565.4]
  wire [7:0] _T_3237; // @[Mux.scala 19:72:@1566.4]
  wire [7:0] _T_3244; // @[Mux.scala 19:72:@1573.4]
  wire [7:0] _T_3246; // @[Mux.scala 19:72:@1574.4]
  wire [7:0] _T_3253; // @[Mux.scala 19:72:@1581.4]
  wire [7:0] _T_3255; // @[Mux.scala 19:72:@1582.4]
  wire [7:0] _T_3262; // @[Mux.scala 19:72:@1589.4]
  wire [7:0] _T_3264; // @[Mux.scala 19:72:@1590.4]
  wire [7:0] _T_3271; // @[Mux.scala 19:72:@1597.4]
  wire [7:0] _T_3273; // @[Mux.scala 19:72:@1598.4]
  wire [7:0] _T_3280; // @[Mux.scala 19:72:@1605.4]
  wire [7:0] _T_3282; // @[Mux.scala 19:72:@1606.4]
  wire [7:0] _T_3289; // @[Mux.scala 19:72:@1613.4]
  wire [7:0] _T_3291; // @[Mux.scala 19:72:@1614.4]
  wire [7:0] _T_3298; // @[Mux.scala 19:72:@1621.4]
  wire [7:0] _T_3300; // @[Mux.scala 19:72:@1622.4]
  wire [7:0] _T_3301; // @[Mux.scala 19:72:@1623.4]
  wire [7:0] _T_3302; // @[Mux.scala 19:72:@1624.4]
  wire [7:0] _T_3303; // @[Mux.scala 19:72:@1625.4]
  wire [7:0] _T_3304; // @[Mux.scala 19:72:@1626.4]
  wire [7:0] _T_3305; // @[Mux.scala 19:72:@1627.4]
  wire [7:0] _T_3306; // @[Mux.scala 19:72:@1628.4]
  wire [7:0] _T_3307; // @[Mux.scala 19:72:@1629.4]
  wire  inputDataPriorityPorts_0_0; // @[Mux.scala 19:72:@1633.4]
  wire  inputDataPriorityPorts_0_1; // @[Mux.scala 19:72:@1635.4]
  wire  inputDataPriorityPorts_0_2; // @[Mux.scala 19:72:@1637.4]
  wire  inputDataPriorityPorts_0_3; // @[Mux.scala 19:72:@1639.4]
  wire  inputDataPriorityPorts_0_4; // @[Mux.scala 19:72:@1641.4]
  wire  inputDataPriorityPorts_0_5; // @[Mux.scala 19:72:@1643.4]
  wire  inputDataPriorityPorts_0_6; // @[Mux.scala 19:72:@1645.4]
  wire  inputDataPriorityPorts_0_7; // @[Mux.scala 19:72:@1647.4]
  wire  _T_3389; // @[StoreQueue.scala 209:52:@1663.6]
  wire  _T_3390; // @[StoreQueue.scala 209:81:@1664.6]
  wire [31:0] _GEN_304; // @[StoreQueue.scala 210:40:@1668.6]
  wire  _GEN_305; // @[StoreQueue.scala 210:40:@1668.6]
  wire  _T_3406; // @[StoreQueue.scala 215:52:@1673.6]
  wire  _T_3407; // @[StoreQueue.scala 215:81:@1674.6]
  wire [31:0] _GEN_306; // @[StoreQueue.scala 216:40:@1678.6]
  wire  _GEN_307; // @[StoreQueue.scala 216:40:@1678.6]
  wire  _GEN_308; // @[StoreQueue.scala 204:35:@1657.4]
  wire  _GEN_309; // @[StoreQueue.scala 204:35:@1657.4]
  wire [31:0] _GEN_310; // @[StoreQueue.scala 204:35:@1657.4]
  wire [31:0] _GEN_311; // @[StoreQueue.scala 204:35:@1657.4]
  wire  _T_3425; // @[StoreQueue.scala 209:52:@1689.6]
  wire  _T_3426; // @[StoreQueue.scala 209:81:@1690.6]
  wire [31:0] _GEN_312; // @[StoreQueue.scala 210:40:@1694.6]
  wire  _GEN_313; // @[StoreQueue.scala 210:40:@1694.6]
  wire  _T_3442; // @[StoreQueue.scala 215:52:@1699.6]
  wire  _T_3443; // @[StoreQueue.scala 215:81:@1700.6]
  wire [31:0] _GEN_314; // @[StoreQueue.scala 216:40:@1704.6]
  wire  _GEN_315; // @[StoreQueue.scala 216:40:@1704.6]
  wire  _GEN_316; // @[StoreQueue.scala 204:35:@1683.4]
  wire  _GEN_317; // @[StoreQueue.scala 204:35:@1683.4]
  wire [31:0] _GEN_318; // @[StoreQueue.scala 204:35:@1683.4]
  wire [31:0] _GEN_319; // @[StoreQueue.scala 204:35:@1683.4]
  wire  _T_3461; // @[StoreQueue.scala 209:52:@1715.6]
  wire  _T_3462; // @[StoreQueue.scala 209:81:@1716.6]
  wire [31:0] _GEN_320; // @[StoreQueue.scala 210:40:@1720.6]
  wire  _GEN_321; // @[StoreQueue.scala 210:40:@1720.6]
  wire  _T_3478; // @[StoreQueue.scala 215:52:@1725.6]
  wire  _T_3479; // @[StoreQueue.scala 215:81:@1726.6]
  wire [31:0] _GEN_322; // @[StoreQueue.scala 216:40:@1730.6]
  wire  _GEN_323; // @[StoreQueue.scala 216:40:@1730.6]
  wire  _GEN_324; // @[StoreQueue.scala 204:35:@1709.4]
  wire  _GEN_325; // @[StoreQueue.scala 204:35:@1709.4]
  wire [31:0] _GEN_326; // @[StoreQueue.scala 204:35:@1709.4]
  wire [31:0] _GEN_327; // @[StoreQueue.scala 204:35:@1709.4]
  wire  _T_3497; // @[StoreQueue.scala 209:52:@1741.6]
  wire  _T_3498; // @[StoreQueue.scala 209:81:@1742.6]
  wire [31:0] _GEN_328; // @[StoreQueue.scala 210:40:@1746.6]
  wire  _GEN_329; // @[StoreQueue.scala 210:40:@1746.6]
  wire  _T_3514; // @[StoreQueue.scala 215:52:@1751.6]
  wire  _T_3515; // @[StoreQueue.scala 215:81:@1752.6]
  wire [31:0] _GEN_330; // @[StoreQueue.scala 216:40:@1756.6]
  wire  _GEN_331; // @[StoreQueue.scala 216:40:@1756.6]
  wire  _GEN_332; // @[StoreQueue.scala 204:35:@1735.4]
  wire  _GEN_333; // @[StoreQueue.scala 204:35:@1735.4]
  wire [31:0] _GEN_334; // @[StoreQueue.scala 204:35:@1735.4]
  wire [31:0] _GEN_335; // @[StoreQueue.scala 204:35:@1735.4]
  wire  _T_3533; // @[StoreQueue.scala 209:52:@1767.6]
  wire  _T_3534; // @[StoreQueue.scala 209:81:@1768.6]
  wire [31:0] _GEN_336; // @[StoreQueue.scala 210:40:@1772.6]
  wire  _GEN_337; // @[StoreQueue.scala 210:40:@1772.6]
  wire  _T_3550; // @[StoreQueue.scala 215:52:@1777.6]
  wire  _T_3551; // @[StoreQueue.scala 215:81:@1778.6]
  wire [31:0] _GEN_338; // @[StoreQueue.scala 216:40:@1782.6]
  wire  _GEN_339; // @[StoreQueue.scala 216:40:@1782.6]
  wire  _GEN_340; // @[StoreQueue.scala 204:35:@1761.4]
  wire  _GEN_341; // @[StoreQueue.scala 204:35:@1761.4]
  wire [31:0] _GEN_342; // @[StoreQueue.scala 204:35:@1761.4]
  wire [31:0] _GEN_343; // @[StoreQueue.scala 204:35:@1761.4]
  wire  _T_3569; // @[StoreQueue.scala 209:52:@1793.6]
  wire  _T_3570; // @[StoreQueue.scala 209:81:@1794.6]
  wire [31:0] _GEN_344; // @[StoreQueue.scala 210:40:@1798.6]
  wire  _GEN_345; // @[StoreQueue.scala 210:40:@1798.6]
  wire  _T_3586; // @[StoreQueue.scala 215:52:@1803.6]
  wire  _T_3587; // @[StoreQueue.scala 215:81:@1804.6]
  wire [31:0] _GEN_346; // @[StoreQueue.scala 216:40:@1808.6]
  wire  _GEN_347; // @[StoreQueue.scala 216:40:@1808.6]
  wire  _GEN_348; // @[StoreQueue.scala 204:35:@1787.4]
  wire  _GEN_349; // @[StoreQueue.scala 204:35:@1787.4]
  wire [31:0] _GEN_350; // @[StoreQueue.scala 204:35:@1787.4]
  wire [31:0] _GEN_351; // @[StoreQueue.scala 204:35:@1787.4]
  wire  _T_3605; // @[StoreQueue.scala 209:52:@1819.6]
  wire  _T_3606; // @[StoreQueue.scala 209:81:@1820.6]
  wire [31:0] _GEN_352; // @[StoreQueue.scala 210:40:@1824.6]
  wire  _GEN_353; // @[StoreQueue.scala 210:40:@1824.6]
  wire  _T_3622; // @[StoreQueue.scala 215:52:@1829.6]
  wire  _T_3623; // @[StoreQueue.scala 215:81:@1830.6]
  wire [31:0] _GEN_354; // @[StoreQueue.scala 216:40:@1834.6]
  wire  _GEN_355; // @[StoreQueue.scala 216:40:@1834.6]
  wire  _GEN_356; // @[StoreQueue.scala 204:35:@1813.4]
  wire  _GEN_357; // @[StoreQueue.scala 204:35:@1813.4]
  wire [31:0] _GEN_358; // @[StoreQueue.scala 204:35:@1813.4]
  wire [31:0] _GEN_359; // @[StoreQueue.scala 204:35:@1813.4]
  wire  _T_3641; // @[StoreQueue.scala 209:52:@1845.6]
  wire  _T_3642; // @[StoreQueue.scala 209:81:@1846.6]
  wire [31:0] _GEN_360; // @[StoreQueue.scala 210:40:@1850.6]
  wire  _GEN_361; // @[StoreQueue.scala 210:40:@1850.6]
  wire  _T_3658; // @[StoreQueue.scala 215:52:@1855.6]
  wire  _T_3659; // @[StoreQueue.scala 215:81:@1856.6]
  wire [31:0] _GEN_362; // @[StoreQueue.scala 216:40:@1860.6]
  wire  _GEN_363; // @[StoreQueue.scala 216:40:@1860.6]
  wire  _GEN_364; // @[StoreQueue.scala 204:35:@1839.4]
  wire  _GEN_365; // @[StoreQueue.scala 204:35:@1839.4]
  wire [31:0] _GEN_366; // @[StoreQueue.scala 204:35:@1839.4]
  wire [31:0] _GEN_367; // @[StoreQueue.scala 204:35:@1839.4]
  wire  _T_3673; // @[StoreQueue.scala 229:23:@1865.4]
  wire [3:0] _T_3676; // @[util.scala 10:8:@1867.6]
  wire [3:0] _GEN_32; // @[util.scala 10:14:@1868.6]
  wire [3:0] _T_3677; // @[util.scala 10:14:@1868.6]
  wire [3:0] _GEN_368; // @[StoreQueue.scala 229:50:@1866.4]
  wire [3:0] _T_3679; // @[util.scala 10:8:@1872.6]
  wire [3:0] _GEN_33; // @[util.scala 10:14:@1873.6]
  wire [3:0] _T_3680; // @[util.scala 10:14:@1873.6]
  wire [3:0] _GEN_369; // @[StoreQueue.scala 233:20:@1871.4]
  wire  _T_3682; // @[StoreQueue.scala 237:84:@1876.4]
  wire  _T_3683; // @[StoreQueue.scala 237:81:@1877.4]
  wire  _T_3685; // @[StoreQueue.scala 237:84:@1878.4]
  wire  _T_3686; // @[StoreQueue.scala 237:81:@1879.4]
  wire  _T_3688; // @[StoreQueue.scala 237:84:@1880.4]
  wire  _T_3689; // @[StoreQueue.scala 237:81:@1881.4]
  wire  _T_3691; // @[StoreQueue.scala 237:84:@1882.4]
  wire  _T_3692; // @[StoreQueue.scala 237:81:@1883.4]
  wire  _T_3694; // @[StoreQueue.scala 237:84:@1884.4]
  wire  _T_3695; // @[StoreQueue.scala 237:81:@1885.4]
  wire  _T_3697; // @[StoreQueue.scala 237:84:@1886.4]
  wire  _T_3698; // @[StoreQueue.scala 237:81:@1887.4]
  wire  _T_3700; // @[StoreQueue.scala 237:84:@1888.4]
  wire  _T_3701; // @[StoreQueue.scala 237:81:@1889.4]
  wire  _T_3703; // @[StoreQueue.scala 237:84:@1890.4]
  wire  _T_3704; // @[StoreQueue.scala 237:81:@1891.4]
  wire  _T_3721; // @[StoreQueue.scala 237:98:@1902.4]
  wire  _T_3722; // @[StoreQueue.scala 237:98:@1903.4]
  wire  _T_3723; // @[StoreQueue.scala 237:98:@1904.4]
  wire  _T_3724; // @[StoreQueue.scala 237:98:@1905.4]
  wire  _T_3725; // @[StoreQueue.scala 237:98:@1906.4]
  wire  _T_3726; // @[StoreQueue.scala 237:98:@1907.4]
  wire [31:0] _GEN_371; // @[StoreQueue.scala 252:21:@1945.4]
  wire [31:0] _GEN_372; // @[StoreQueue.scala 252:21:@1945.4]
  wire [31:0] _GEN_373; // @[StoreQueue.scala 252:21:@1945.4]
  wire [31:0] _GEN_374; // @[StoreQueue.scala 252:21:@1945.4]
  wire [31:0] _GEN_375; // @[StoreQueue.scala 252:21:@1945.4]
  wire [31:0] _GEN_376; // @[StoreQueue.scala 252:21:@1945.4]
  assign _GEN_378 = {{2'd0}, tail}; // @[util.scala 14:20:@101.4]
  assign _T_948 = 5'h8 - _GEN_378; // @[util.scala 14:20:@101.4]
  assign _T_949 = $unsigned(_T_948); // @[util.scala 14:20:@102.4]
  assign _T_950 = _T_949[4:0]; // @[util.scala 14:20:@103.4]
  assign _GEN_0 = _T_950 % 5'h8; // @[util.scala 14:25:@104.4]
  assign _T_951 = _GEN_0[3:0]; // @[util.scala 14:25:@104.4]
  assign _GEN_379 = {{1'd0}, io_bbNumStores}; // @[StoreQueue.scala 70:46:@105.4]
  assign _T_952 = _T_951 < _GEN_379; // @[StoreQueue.scala 70:46:@105.4]
  assign initBits_0 = _T_952 & io_bbStart; // @[StoreQueue.scala 70:64:@106.4]
  assign _T_957 = 5'h9 - _GEN_378; // @[util.scala 14:20:@108.4]
  assign _T_958 = $unsigned(_T_957); // @[util.scala 14:20:@109.4]
  assign _T_959 = _T_958[4:0]; // @[util.scala 14:20:@110.4]
  assign _GEN_8 = _T_959 % 5'h8; // @[util.scala 14:25:@111.4]
  assign _T_960 = _GEN_8[3:0]; // @[util.scala 14:25:@111.4]
  assign _T_961 = _T_960 < _GEN_379; // @[StoreQueue.scala 70:46:@112.4]
  assign initBits_1 = _T_961 & io_bbStart; // @[StoreQueue.scala 70:64:@113.4]
  assign _T_966 = 5'ha - _GEN_378; // @[util.scala 14:20:@115.4]
  assign _T_967 = $unsigned(_T_966); // @[util.scala 14:20:@116.4]
  assign _T_968 = _T_967[4:0]; // @[util.scala 14:20:@117.4]
  assign _GEN_9 = _T_968 % 5'h8; // @[util.scala 14:25:@118.4]
  assign _T_969 = _GEN_9[3:0]; // @[util.scala 14:25:@118.4]
  assign _T_970 = _T_969 < _GEN_379; // @[StoreQueue.scala 70:46:@119.4]
  assign initBits_2 = _T_970 & io_bbStart; // @[StoreQueue.scala 70:64:@120.4]
  assign _T_975 = 5'hb - _GEN_378; // @[util.scala 14:20:@122.4]
  assign _T_976 = $unsigned(_T_975); // @[util.scala 14:20:@123.4]
  assign _T_977 = _T_976[4:0]; // @[util.scala 14:20:@124.4]
  assign _GEN_10 = _T_977 % 5'h8; // @[util.scala 14:25:@125.4]
  assign _T_978 = _GEN_10[3:0]; // @[util.scala 14:25:@125.4]
  assign _T_979 = _T_978 < _GEN_379; // @[StoreQueue.scala 70:46:@126.4]
  assign initBits_3 = _T_979 & io_bbStart; // @[StoreQueue.scala 70:64:@127.4]
  assign _T_984 = 5'hc - _GEN_378; // @[util.scala 14:20:@129.4]
  assign _T_985 = $unsigned(_T_984); // @[util.scala 14:20:@130.4]
  assign _T_986 = _T_985[4:0]; // @[util.scala 14:20:@131.4]
  assign _GEN_11 = _T_986 % 5'h8; // @[util.scala 14:25:@132.4]
  assign _T_987 = _GEN_11[3:0]; // @[util.scala 14:25:@132.4]
  assign _T_988 = _T_987 < _GEN_379; // @[StoreQueue.scala 70:46:@133.4]
  assign initBits_4 = _T_988 & io_bbStart; // @[StoreQueue.scala 70:64:@134.4]
  assign _T_993 = 5'hd - _GEN_378; // @[util.scala 14:20:@136.4]
  assign _T_994 = $unsigned(_T_993); // @[util.scala 14:20:@137.4]
  assign _T_995 = _T_994[4:0]; // @[util.scala 14:20:@138.4]
  assign _GEN_12 = _T_995 % 5'h8; // @[util.scala 14:25:@139.4]
  assign _T_996 = _GEN_12[3:0]; // @[util.scala 14:25:@139.4]
  assign _T_997 = _T_996 < _GEN_379; // @[StoreQueue.scala 70:46:@140.4]
  assign initBits_5 = _T_997 & io_bbStart; // @[StoreQueue.scala 70:64:@141.4]
  assign _T_1002 = 5'he - _GEN_378; // @[util.scala 14:20:@143.4]
  assign _T_1003 = $unsigned(_T_1002); // @[util.scala 14:20:@144.4]
  assign _T_1004 = _T_1003[4:0]; // @[util.scala 14:20:@145.4]
  assign _GEN_13 = _T_1004 % 5'h8; // @[util.scala 14:25:@146.4]
  assign _T_1005 = _GEN_13[3:0]; // @[util.scala 14:25:@146.4]
  assign _T_1006 = _T_1005 < _GEN_379; // @[StoreQueue.scala 70:46:@147.4]
  assign initBits_6 = _T_1006 & io_bbStart; // @[StoreQueue.scala 70:64:@148.4]
  assign _T_1011 = 5'hf - _GEN_378; // @[util.scala 14:20:@150.4]
  assign _T_1012 = $unsigned(_T_1011); // @[util.scala 14:20:@151.4]
  assign _T_1013 = _T_1012[4:0]; // @[util.scala 14:20:@152.4]
  assign _GEN_14 = _T_1013 % 5'h8; // @[util.scala 14:25:@153.4]
  assign _T_1014 = _GEN_14[3:0]; // @[util.scala 14:25:@153.4]
  assign _T_1015 = _T_1014 < _GEN_379; // @[StoreQueue.scala 70:46:@154.4]
  assign initBits_7 = _T_1015 & io_bbStart; // @[StoreQueue.scala 70:64:@155.4]
  assign _T_1030 = allocatedEntries_0 | initBits_0; // @[StoreQueue.scala 72:78:@165.4]
  assign _T_1031 = allocatedEntries_1 | initBits_1; // @[StoreQueue.scala 72:78:@166.4]
  assign _T_1032 = allocatedEntries_2 | initBits_2; // @[StoreQueue.scala 72:78:@167.4]
  assign _T_1033 = allocatedEntries_3 | initBits_3; // @[StoreQueue.scala 72:78:@168.4]
  assign _T_1034 = allocatedEntries_4 | initBits_4; // @[StoreQueue.scala 72:78:@169.4]
  assign _T_1035 = allocatedEntries_5 | initBits_5; // @[StoreQueue.scala 72:78:@170.4]
  assign _T_1036 = allocatedEntries_6 | initBits_6; // @[StoreQueue.scala 72:78:@171.4]
  assign _T_1037 = allocatedEntries_7 | initBits_7; // @[StoreQueue.scala 72:78:@172.4]
  assign _T_1060 = _T_951[2:0]; // @[:@196.6]
  assign _GEN_1 = 3'h1 == _T_1060 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_2 = 3'h2 == _T_1060 ? io_bbStoreOffsets_2 : _GEN_1; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_3 = 3'h3 == _T_1060 ? io_bbStoreOffsets_3 : _GEN_2; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_4 = 3'h4 == _T_1060 ? io_bbStoreOffsets_4 : _GEN_3; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_5 = 3'h5 == _T_1060 ? io_bbStoreOffsets_5 : _GEN_4; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_6 = 3'h6 == _T_1060 ? io_bbStoreOffsets_6 : _GEN_5; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_7 = 3'h7 == _T_1060 ? io_bbStoreOffsets_7 : _GEN_6; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_16 = initBits_0 ? _GEN_7 : offsetQ_0; // @[StoreQueue.scala 75:25:@190.4]
  assign _GEN_17 = initBits_0 ? 1'h0 : portQ_0; // @[StoreQueue.scala 75:25:@190.4]
  assign _T_1078 = _T_960[2:0]; // @[:@212.6]
  assign _GEN_19 = 3'h1 == _T_1078 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_20 = 3'h2 == _T_1078 ? io_bbStoreOffsets_2 : _GEN_19; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_21 = 3'h3 == _T_1078 ? io_bbStoreOffsets_3 : _GEN_20; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_22 = 3'h4 == _T_1078 ? io_bbStoreOffsets_4 : _GEN_21; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_23 = 3'h5 == _T_1078 ? io_bbStoreOffsets_5 : _GEN_22; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_24 = 3'h6 == _T_1078 ? io_bbStoreOffsets_6 : _GEN_23; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_25 = 3'h7 == _T_1078 ? io_bbStoreOffsets_7 : _GEN_24; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_34 = initBits_1 ? _GEN_25 : offsetQ_1; // @[StoreQueue.scala 75:25:@206.4]
  assign _GEN_35 = initBits_1 ? 1'h0 : portQ_1; // @[StoreQueue.scala 75:25:@206.4]
  assign _T_1096 = _T_969[2:0]; // @[:@228.6]
  assign _GEN_37 = 3'h1 == _T_1096 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_38 = 3'h2 == _T_1096 ? io_bbStoreOffsets_2 : _GEN_37; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_39 = 3'h3 == _T_1096 ? io_bbStoreOffsets_3 : _GEN_38; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_40 = 3'h4 == _T_1096 ? io_bbStoreOffsets_4 : _GEN_39; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_41 = 3'h5 == _T_1096 ? io_bbStoreOffsets_5 : _GEN_40; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_42 = 3'h6 == _T_1096 ? io_bbStoreOffsets_6 : _GEN_41; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_43 = 3'h7 == _T_1096 ? io_bbStoreOffsets_7 : _GEN_42; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_52 = initBits_2 ? _GEN_43 : offsetQ_2; // @[StoreQueue.scala 75:25:@222.4]
  assign _GEN_53 = initBits_2 ? 1'h0 : portQ_2; // @[StoreQueue.scala 75:25:@222.4]
  assign _T_1114 = _T_978[2:0]; // @[:@244.6]
  assign _GEN_55 = 3'h1 == _T_1114 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_56 = 3'h2 == _T_1114 ? io_bbStoreOffsets_2 : _GEN_55; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_57 = 3'h3 == _T_1114 ? io_bbStoreOffsets_3 : _GEN_56; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_58 = 3'h4 == _T_1114 ? io_bbStoreOffsets_4 : _GEN_57; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_59 = 3'h5 == _T_1114 ? io_bbStoreOffsets_5 : _GEN_58; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_60 = 3'h6 == _T_1114 ? io_bbStoreOffsets_6 : _GEN_59; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_61 = 3'h7 == _T_1114 ? io_bbStoreOffsets_7 : _GEN_60; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_70 = initBits_3 ? _GEN_61 : offsetQ_3; // @[StoreQueue.scala 75:25:@238.4]
  assign _GEN_71 = initBits_3 ? 1'h0 : portQ_3; // @[StoreQueue.scala 75:25:@238.4]
  assign _T_1132 = _T_987[2:0]; // @[:@260.6]
  assign _GEN_73 = 3'h1 == _T_1132 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_74 = 3'h2 == _T_1132 ? io_bbStoreOffsets_2 : _GEN_73; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_75 = 3'h3 == _T_1132 ? io_bbStoreOffsets_3 : _GEN_74; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_76 = 3'h4 == _T_1132 ? io_bbStoreOffsets_4 : _GEN_75; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_77 = 3'h5 == _T_1132 ? io_bbStoreOffsets_5 : _GEN_76; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_78 = 3'h6 == _T_1132 ? io_bbStoreOffsets_6 : _GEN_77; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_79 = 3'h7 == _T_1132 ? io_bbStoreOffsets_7 : _GEN_78; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_88 = initBits_4 ? _GEN_79 : offsetQ_4; // @[StoreQueue.scala 75:25:@254.4]
  assign _GEN_89 = initBits_4 ? 1'h0 : portQ_4; // @[StoreQueue.scala 75:25:@254.4]
  assign _T_1150 = _T_996[2:0]; // @[:@276.6]
  assign _GEN_91 = 3'h1 == _T_1150 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_92 = 3'h2 == _T_1150 ? io_bbStoreOffsets_2 : _GEN_91; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_93 = 3'h3 == _T_1150 ? io_bbStoreOffsets_3 : _GEN_92; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_94 = 3'h4 == _T_1150 ? io_bbStoreOffsets_4 : _GEN_93; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_95 = 3'h5 == _T_1150 ? io_bbStoreOffsets_5 : _GEN_94; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_96 = 3'h6 == _T_1150 ? io_bbStoreOffsets_6 : _GEN_95; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_97 = 3'h7 == _T_1150 ? io_bbStoreOffsets_7 : _GEN_96; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_106 = initBits_5 ? _GEN_97 : offsetQ_5; // @[StoreQueue.scala 75:25:@270.4]
  assign _GEN_107 = initBits_5 ? 1'h0 : portQ_5; // @[StoreQueue.scala 75:25:@270.4]
  assign _T_1168 = _T_1005[2:0]; // @[:@292.6]
  assign _GEN_109 = 3'h1 == _T_1168 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_110 = 3'h2 == _T_1168 ? io_bbStoreOffsets_2 : _GEN_109; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_111 = 3'h3 == _T_1168 ? io_bbStoreOffsets_3 : _GEN_110; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_112 = 3'h4 == _T_1168 ? io_bbStoreOffsets_4 : _GEN_111; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_113 = 3'h5 == _T_1168 ? io_bbStoreOffsets_5 : _GEN_112; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_114 = 3'h6 == _T_1168 ? io_bbStoreOffsets_6 : _GEN_113; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_115 = 3'h7 == _T_1168 ? io_bbStoreOffsets_7 : _GEN_114; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_124 = initBits_6 ? _GEN_115 : offsetQ_6; // @[StoreQueue.scala 75:25:@286.4]
  assign _GEN_125 = initBits_6 ? 1'h0 : portQ_6; // @[StoreQueue.scala 75:25:@286.4]
  assign _T_1186 = _T_1014[2:0]; // @[:@308.6]
  assign _GEN_127 = 3'h1 == _T_1186 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_128 = 3'h2 == _T_1186 ? io_bbStoreOffsets_2 : _GEN_127; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_129 = 3'h3 == _T_1186 ? io_bbStoreOffsets_3 : _GEN_128; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_130 = 3'h4 == _T_1186 ? io_bbStoreOffsets_4 : _GEN_129; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_131 = 3'h5 == _T_1186 ? io_bbStoreOffsets_5 : _GEN_130; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_132 = 3'h6 == _T_1186 ? io_bbStoreOffsets_6 : _GEN_131; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_133 = 3'h7 == _T_1186 ? io_bbStoreOffsets_7 : _GEN_132; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_142 = initBits_7 ? _GEN_133 : offsetQ_7; // @[StoreQueue.scala 75:25:@302.4]
  assign _GEN_143 = initBits_7 ? 1'h0 : portQ_7; // @[StoreQueue.scala 75:25:@302.4]
  assign _T_1208 = _GEN_7 + 3'h1; // @[util.scala 10:8:@327.6]
  assign _GEN_15 = _T_1208 % 4'h8; // @[util.scala 10:14:@328.6]
  assign _T_1209 = _GEN_15[3:0]; // @[util.scala 10:14:@328.6]
  assign _GEN_411 = {{1'd0}, io_loadTail}; // @[StoreQueue.scala 96:56:@329.6]
  assign _T_1210 = _T_1209 == _GEN_411; // @[StoreQueue.scala 96:56:@329.6]
  assign _T_1211 = io_loadEmpty & _T_1210; // @[StoreQueue.scala 95:50:@330.6]
  assign _T_1213 = _T_1211 == 1'h0; // @[StoreQueue.scala 95:35:@331.6]
  assign _T_1215 = previousLoadHead <= offsetQ_0; // @[StoreQueue.scala 100:35:@339.8]
  assign _T_1216 = offsetQ_0 < io_loadHead; // @[StoreQueue.scala 100:87:@340.8]
  assign _T_1217 = _T_1215 & _T_1216; // @[StoreQueue.scala 100:61:@341.8]
  assign _T_1219 = previousLoadHead > io_loadHead; // @[StoreQueue.scala 102:35:@346.10]
  assign _T_1220 = io_loadHead <= offsetQ_0; // @[StoreQueue.scala 103:23:@347.10]
  assign _T_1221 = offsetQ_0 < previousLoadHead; // @[StoreQueue.scala 103:75:@348.10]
  assign _T_1222 = _T_1220 & _T_1221; // @[StoreQueue.scala 103:49:@349.10]
  assign _T_1224 = _T_1222 == 1'h0; // @[StoreQueue.scala 103:9:@350.10]
  assign _T_1225 = _T_1219 & _T_1224; // @[StoreQueue.scala 102:49:@351.10]
  assign _GEN_152 = _T_1225 ? 1'h0 : checkBits_0; // @[StoreQueue.scala 103:96:@352.10]
  assign _GEN_153 = _T_1217 ? 1'h0 : _GEN_152; // @[StoreQueue.scala 100:102:@342.8]
  assign _GEN_154 = io_loadEmpty ? 1'h0 : _GEN_153; // @[StoreQueue.scala 98:26:@335.6]
  assign _GEN_155 = initBits_0 ? _T_1213 : _GEN_154; // @[StoreQueue.scala 94:35:@320.4]
  assign _T_1238 = _GEN_25 + 3'h1; // @[util.scala 10:8:@363.6]
  assign _GEN_18 = _T_1238 % 4'h8; // @[util.scala 10:14:@364.6]
  assign _T_1239 = _GEN_18[3:0]; // @[util.scala 10:14:@364.6]
  assign _T_1240 = _T_1239 == _GEN_411; // @[StoreQueue.scala 96:56:@365.6]
  assign _T_1241 = io_loadEmpty & _T_1240; // @[StoreQueue.scala 95:50:@366.6]
  assign _T_1243 = _T_1241 == 1'h0; // @[StoreQueue.scala 95:35:@367.6]
  assign _T_1245 = previousLoadHead <= offsetQ_1; // @[StoreQueue.scala 100:35:@375.8]
  assign _T_1246 = offsetQ_1 < io_loadHead; // @[StoreQueue.scala 100:87:@376.8]
  assign _T_1247 = _T_1245 & _T_1246; // @[StoreQueue.scala 100:61:@377.8]
  assign _T_1250 = io_loadHead <= offsetQ_1; // @[StoreQueue.scala 103:23:@383.10]
  assign _T_1251 = offsetQ_1 < previousLoadHead; // @[StoreQueue.scala 103:75:@384.10]
  assign _T_1252 = _T_1250 & _T_1251; // @[StoreQueue.scala 103:49:@385.10]
  assign _T_1254 = _T_1252 == 1'h0; // @[StoreQueue.scala 103:9:@386.10]
  assign _T_1255 = _T_1219 & _T_1254; // @[StoreQueue.scala 102:49:@387.10]
  assign _GEN_164 = _T_1255 ? 1'h0 : checkBits_1; // @[StoreQueue.scala 103:96:@388.10]
  assign _GEN_165 = _T_1247 ? 1'h0 : _GEN_164; // @[StoreQueue.scala 100:102:@378.8]
  assign _GEN_166 = io_loadEmpty ? 1'h0 : _GEN_165; // @[StoreQueue.scala 98:26:@371.6]
  assign _GEN_167 = initBits_1 ? _T_1243 : _GEN_166; // @[StoreQueue.scala 94:35:@356.4]
  assign _T_1268 = _GEN_43 + 3'h1; // @[util.scala 10:8:@399.6]
  assign _GEN_26 = _T_1268 % 4'h8; // @[util.scala 10:14:@400.6]
  assign _T_1269 = _GEN_26[3:0]; // @[util.scala 10:14:@400.6]
  assign _T_1270 = _T_1269 == _GEN_411; // @[StoreQueue.scala 96:56:@401.6]
  assign _T_1271 = io_loadEmpty & _T_1270; // @[StoreQueue.scala 95:50:@402.6]
  assign _T_1273 = _T_1271 == 1'h0; // @[StoreQueue.scala 95:35:@403.6]
  assign _T_1275 = previousLoadHead <= offsetQ_2; // @[StoreQueue.scala 100:35:@411.8]
  assign _T_1276 = offsetQ_2 < io_loadHead; // @[StoreQueue.scala 100:87:@412.8]
  assign _T_1277 = _T_1275 & _T_1276; // @[StoreQueue.scala 100:61:@413.8]
  assign _T_1280 = io_loadHead <= offsetQ_2; // @[StoreQueue.scala 103:23:@419.10]
  assign _T_1281 = offsetQ_2 < previousLoadHead; // @[StoreQueue.scala 103:75:@420.10]
  assign _T_1282 = _T_1280 & _T_1281; // @[StoreQueue.scala 103:49:@421.10]
  assign _T_1284 = _T_1282 == 1'h0; // @[StoreQueue.scala 103:9:@422.10]
  assign _T_1285 = _T_1219 & _T_1284; // @[StoreQueue.scala 102:49:@423.10]
  assign _GEN_176 = _T_1285 ? 1'h0 : checkBits_2; // @[StoreQueue.scala 103:96:@424.10]
  assign _GEN_177 = _T_1277 ? 1'h0 : _GEN_176; // @[StoreQueue.scala 100:102:@414.8]
  assign _GEN_178 = io_loadEmpty ? 1'h0 : _GEN_177; // @[StoreQueue.scala 98:26:@407.6]
  assign _GEN_179 = initBits_2 ? _T_1273 : _GEN_178; // @[StoreQueue.scala 94:35:@392.4]
  assign _T_1298 = _GEN_61 + 3'h1; // @[util.scala 10:8:@435.6]
  assign _GEN_27 = _T_1298 % 4'h8; // @[util.scala 10:14:@436.6]
  assign _T_1299 = _GEN_27[3:0]; // @[util.scala 10:14:@436.6]
  assign _T_1300 = _T_1299 == _GEN_411; // @[StoreQueue.scala 96:56:@437.6]
  assign _T_1301 = io_loadEmpty & _T_1300; // @[StoreQueue.scala 95:50:@438.6]
  assign _T_1303 = _T_1301 == 1'h0; // @[StoreQueue.scala 95:35:@439.6]
  assign _T_1305 = previousLoadHead <= offsetQ_3; // @[StoreQueue.scala 100:35:@447.8]
  assign _T_1306 = offsetQ_3 < io_loadHead; // @[StoreQueue.scala 100:87:@448.8]
  assign _T_1307 = _T_1305 & _T_1306; // @[StoreQueue.scala 100:61:@449.8]
  assign _T_1310 = io_loadHead <= offsetQ_3; // @[StoreQueue.scala 103:23:@455.10]
  assign _T_1311 = offsetQ_3 < previousLoadHead; // @[StoreQueue.scala 103:75:@456.10]
  assign _T_1312 = _T_1310 & _T_1311; // @[StoreQueue.scala 103:49:@457.10]
  assign _T_1314 = _T_1312 == 1'h0; // @[StoreQueue.scala 103:9:@458.10]
  assign _T_1315 = _T_1219 & _T_1314; // @[StoreQueue.scala 102:49:@459.10]
  assign _GEN_188 = _T_1315 ? 1'h0 : checkBits_3; // @[StoreQueue.scala 103:96:@460.10]
  assign _GEN_189 = _T_1307 ? 1'h0 : _GEN_188; // @[StoreQueue.scala 100:102:@450.8]
  assign _GEN_190 = io_loadEmpty ? 1'h0 : _GEN_189; // @[StoreQueue.scala 98:26:@443.6]
  assign _GEN_191 = initBits_3 ? _T_1303 : _GEN_190; // @[StoreQueue.scala 94:35:@428.4]
  assign _T_1328 = _GEN_79 + 3'h1; // @[util.scala 10:8:@471.6]
  assign _GEN_28 = _T_1328 % 4'h8; // @[util.scala 10:14:@472.6]
  assign _T_1329 = _GEN_28[3:0]; // @[util.scala 10:14:@472.6]
  assign _T_1330 = _T_1329 == _GEN_411; // @[StoreQueue.scala 96:56:@473.6]
  assign _T_1331 = io_loadEmpty & _T_1330; // @[StoreQueue.scala 95:50:@474.6]
  assign _T_1333 = _T_1331 == 1'h0; // @[StoreQueue.scala 95:35:@475.6]
  assign _T_1335 = previousLoadHead <= offsetQ_4; // @[StoreQueue.scala 100:35:@483.8]
  assign _T_1336 = offsetQ_4 < io_loadHead; // @[StoreQueue.scala 100:87:@484.8]
  assign _T_1337 = _T_1335 & _T_1336; // @[StoreQueue.scala 100:61:@485.8]
  assign _T_1340 = io_loadHead <= offsetQ_4; // @[StoreQueue.scala 103:23:@491.10]
  assign _T_1341 = offsetQ_4 < previousLoadHead; // @[StoreQueue.scala 103:75:@492.10]
  assign _T_1342 = _T_1340 & _T_1341; // @[StoreQueue.scala 103:49:@493.10]
  assign _T_1344 = _T_1342 == 1'h0; // @[StoreQueue.scala 103:9:@494.10]
  assign _T_1345 = _T_1219 & _T_1344; // @[StoreQueue.scala 102:49:@495.10]
  assign _GEN_200 = _T_1345 ? 1'h0 : checkBits_4; // @[StoreQueue.scala 103:96:@496.10]
  assign _GEN_201 = _T_1337 ? 1'h0 : _GEN_200; // @[StoreQueue.scala 100:102:@486.8]
  assign _GEN_202 = io_loadEmpty ? 1'h0 : _GEN_201; // @[StoreQueue.scala 98:26:@479.6]
  assign _GEN_203 = initBits_4 ? _T_1333 : _GEN_202; // @[StoreQueue.scala 94:35:@464.4]
  assign _T_1358 = _GEN_97 + 3'h1; // @[util.scala 10:8:@507.6]
  assign _GEN_29 = _T_1358 % 4'h8; // @[util.scala 10:14:@508.6]
  assign _T_1359 = _GEN_29[3:0]; // @[util.scala 10:14:@508.6]
  assign _T_1360 = _T_1359 == _GEN_411; // @[StoreQueue.scala 96:56:@509.6]
  assign _T_1361 = io_loadEmpty & _T_1360; // @[StoreQueue.scala 95:50:@510.6]
  assign _T_1363 = _T_1361 == 1'h0; // @[StoreQueue.scala 95:35:@511.6]
  assign _T_1365 = previousLoadHead <= offsetQ_5; // @[StoreQueue.scala 100:35:@519.8]
  assign _T_1366 = offsetQ_5 < io_loadHead; // @[StoreQueue.scala 100:87:@520.8]
  assign _T_1367 = _T_1365 & _T_1366; // @[StoreQueue.scala 100:61:@521.8]
  assign _T_1370 = io_loadHead <= offsetQ_5; // @[StoreQueue.scala 103:23:@527.10]
  assign _T_1371 = offsetQ_5 < previousLoadHead; // @[StoreQueue.scala 103:75:@528.10]
  assign _T_1372 = _T_1370 & _T_1371; // @[StoreQueue.scala 103:49:@529.10]
  assign _T_1374 = _T_1372 == 1'h0; // @[StoreQueue.scala 103:9:@530.10]
  assign _T_1375 = _T_1219 & _T_1374; // @[StoreQueue.scala 102:49:@531.10]
  assign _GEN_212 = _T_1375 ? 1'h0 : checkBits_5; // @[StoreQueue.scala 103:96:@532.10]
  assign _GEN_213 = _T_1367 ? 1'h0 : _GEN_212; // @[StoreQueue.scala 100:102:@522.8]
  assign _GEN_214 = io_loadEmpty ? 1'h0 : _GEN_213; // @[StoreQueue.scala 98:26:@515.6]
  assign _GEN_215 = initBits_5 ? _T_1363 : _GEN_214; // @[StoreQueue.scala 94:35:@500.4]
  assign _T_1388 = _GEN_115 + 3'h1; // @[util.scala 10:8:@543.6]
  assign _GEN_30 = _T_1388 % 4'h8; // @[util.scala 10:14:@544.6]
  assign _T_1389 = _GEN_30[3:0]; // @[util.scala 10:14:@544.6]
  assign _T_1390 = _T_1389 == _GEN_411; // @[StoreQueue.scala 96:56:@545.6]
  assign _T_1391 = io_loadEmpty & _T_1390; // @[StoreQueue.scala 95:50:@546.6]
  assign _T_1393 = _T_1391 == 1'h0; // @[StoreQueue.scala 95:35:@547.6]
  assign _T_1395 = previousLoadHead <= offsetQ_6; // @[StoreQueue.scala 100:35:@555.8]
  assign _T_1396 = offsetQ_6 < io_loadHead; // @[StoreQueue.scala 100:87:@556.8]
  assign _T_1397 = _T_1395 & _T_1396; // @[StoreQueue.scala 100:61:@557.8]
  assign _T_1400 = io_loadHead <= offsetQ_6; // @[StoreQueue.scala 103:23:@563.10]
  assign _T_1401 = offsetQ_6 < previousLoadHead; // @[StoreQueue.scala 103:75:@564.10]
  assign _T_1402 = _T_1400 & _T_1401; // @[StoreQueue.scala 103:49:@565.10]
  assign _T_1404 = _T_1402 == 1'h0; // @[StoreQueue.scala 103:9:@566.10]
  assign _T_1405 = _T_1219 & _T_1404; // @[StoreQueue.scala 102:49:@567.10]
  assign _GEN_224 = _T_1405 ? 1'h0 : checkBits_6; // @[StoreQueue.scala 103:96:@568.10]
  assign _GEN_225 = _T_1397 ? 1'h0 : _GEN_224; // @[StoreQueue.scala 100:102:@558.8]
  assign _GEN_226 = io_loadEmpty ? 1'h0 : _GEN_225; // @[StoreQueue.scala 98:26:@551.6]
  assign _GEN_227 = initBits_6 ? _T_1393 : _GEN_226; // @[StoreQueue.scala 94:35:@536.4]
  assign _T_1418 = _GEN_133 + 3'h1; // @[util.scala 10:8:@579.6]
  assign _GEN_31 = _T_1418 % 4'h8; // @[util.scala 10:14:@580.6]
  assign _T_1419 = _GEN_31[3:0]; // @[util.scala 10:14:@580.6]
  assign _T_1420 = _T_1419 == _GEN_411; // @[StoreQueue.scala 96:56:@581.6]
  assign _T_1421 = io_loadEmpty & _T_1420; // @[StoreQueue.scala 95:50:@582.6]
  assign _T_1423 = _T_1421 == 1'h0; // @[StoreQueue.scala 95:35:@583.6]
  assign _T_1425 = previousLoadHead <= offsetQ_7; // @[StoreQueue.scala 100:35:@591.8]
  assign _T_1426 = offsetQ_7 < io_loadHead; // @[StoreQueue.scala 100:87:@592.8]
  assign _T_1427 = _T_1425 & _T_1426; // @[StoreQueue.scala 100:61:@593.8]
  assign _T_1430 = io_loadHead <= offsetQ_7; // @[StoreQueue.scala 103:23:@599.10]
  assign _T_1431 = offsetQ_7 < previousLoadHead; // @[StoreQueue.scala 103:75:@600.10]
  assign _T_1432 = _T_1430 & _T_1431; // @[StoreQueue.scala 103:49:@601.10]
  assign _T_1434 = _T_1432 == 1'h0; // @[StoreQueue.scala 103:9:@602.10]
  assign _T_1435 = _T_1219 & _T_1434; // @[StoreQueue.scala 102:49:@603.10]
  assign _GEN_236 = _T_1435 ? 1'h0 : checkBits_7; // @[StoreQueue.scala 103:96:@604.10]
  assign _GEN_237 = _T_1427 ? 1'h0 : _GEN_236; // @[StoreQueue.scala 100:102:@594.8]
  assign _GEN_238 = io_loadEmpty ? 1'h0 : _GEN_237; // @[StoreQueue.scala 98:26:@587.6]
  assign _GEN_239 = initBits_7 ? _T_1423 : _GEN_238; // @[StoreQueue.scala 94:35:@572.4]
  assign _T_1437 = io_loadHead < io_loadTail; // @[StoreQueue.scala 119:103:@608.4]
  assign _T_1439 = io_loadHead <= 3'h0; // @[StoreQueue.scala 120:17:@609.4]
  assign _T_1441 = 3'h0 < io_loadTail; // @[StoreQueue.scala 120:35:@610.4]
  assign _T_1442 = _T_1439 & _T_1441; // @[StoreQueue.scala 120:26:@611.4]
  assign _T_1444 = io_loadEmpty == 1'h0; // @[StoreQueue.scala 120:50:@612.4]
  assign _T_1446 = io_loadTail <= 3'h0; // @[StoreQueue.scala 120:81:@613.4]
  assign _T_1448 = 3'h0 < io_loadHead; // @[StoreQueue.scala 120:99:@614.4]
  assign _T_1449 = _T_1446 & _T_1448; // @[StoreQueue.scala 120:90:@615.4]
  assign _T_1451 = _T_1449 == 1'h0; // @[StoreQueue.scala 120:67:@616.4]
  assign _T_1452 = _T_1444 & _T_1451; // @[StoreQueue.scala 120:64:@617.4]
  assign validEntriesInLoadQ_0 = _T_1437 ? _T_1442 : _T_1452; // @[StoreQueue.scala 119:90:@618.4]
  assign _T_1456 = io_loadHead <= 3'h1; // @[StoreQueue.scala 120:17:@620.4]
  assign _T_1458 = 3'h1 < io_loadTail; // @[StoreQueue.scala 120:35:@621.4]
  assign _T_1459 = _T_1456 & _T_1458; // @[StoreQueue.scala 120:26:@622.4]
  assign _T_1463 = io_loadTail <= 3'h1; // @[StoreQueue.scala 120:81:@624.4]
  assign _T_1465 = 3'h1 < io_loadHead; // @[StoreQueue.scala 120:99:@625.4]
  assign _T_1466 = _T_1463 & _T_1465; // @[StoreQueue.scala 120:90:@626.4]
  assign _T_1468 = _T_1466 == 1'h0; // @[StoreQueue.scala 120:67:@627.4]
  assign _T_1469 = _T_1444 & _T_1468; // @[StoreQueue.scala 120:64:@628.4]
  assign validEntriesInLoadQ_1 = _T_1437 ? _T_1459 : _T_1469; // @[StoreQueue.scala 119:90:@629.4]
  assign _T_1473 = io_loadHead <= 3'h2; // @[StoreQueue.scala 120:17:@631.4]
  assign _T_1475 = 3'h2 < io_loadTail; // @[StoreQueue.scala 120:35:@632.4]
  assign _T_1476 = _T_1473 & _T_1475; // @[StoreQueue.scala 120:26:@633.4]
  assign _T_1480 = io_loadTail <= 3'h2; // @[StoreQueue.scala 120:81:@635.4]
  assign _T_1482 = 3'h2 < io_loadHead; // @[StoreQueue.scala 120:99:@636.4]
  assign _T_1483 = _T_1480 & _T_1482; // @[StoreQueue.scala 120:90:@637.4]
  assign _T_1485 = _T_1483 == 1'h0; // @[StoreQueue.scala 120:67:@638.4]
  assign _T_1486 = _T_1444 & _T_1485; // @[StoreQueue.scala 120:64:@639.4]
  assign validEntriesInLoadQ_2 = _T_1437 ? _T_1476 : _T_1486; // @[StoreQueue.scala 119:90:@640.4]
  assign _T_1490 = io_loadHead <= 3'h3; // @[StoreQueue.scala 120:17:@642.4]
  assign _T_1492 = 3'h3 < io_loadTail; // @[StoreQueue.scala 120:35:@643.4]
  assign _T_1493 = _T_1490 & _T_1492; // @[StoreQueue.scala 120:26:@644.4]
  assign _T_1497 = io_loadTail <= 3'h3; // @[StoreQueue.scala 120:81:@646.4]
  assign _T_1499 = 3'h3 < io_loadHead; // @[StoreQueue.scala 120:99:@647.4]
  assign _T_1500 = _T_1497 & _T_1499; // @[StoreQueue.scala 120:90:@648.4]
  assign _T_1502 = _T_1500 == 1'h0; // @[StoreQueue.scala 120:67:@649.4]
  assign _T_1503 = _T_1444 & _T_1502; // @[StoreQueue.scala 120:64:@650.4]
  assign validEntriesInLoadQ_3 = _T_1437 ? _T_1493 : _T_1503; // @[StoreQueue.scala 119:90:@651.4]
  assign _T_1507 = io_loadHead <= 3'h4; // @[StoreQueue.scala 120:17:@653.4]
  assign _T_1509 = 3'h4 < io_loadTail; // @[StoreQueue.scala 120:35:@654.4]
  assign _T_1510 = _T_1507 & _T_1509; // @[StoreQueue.scala 120:26:@655.4]
  assign _T_1514 = io_loadTail <= 3'h4; // @[StoreQueue.scala 120:81:@657.4]
  assign _T_1516 = 3'h4 < io_loadHead; // @[StoreQueue.scala 120:99:@658.4]
  assign _T_1517 = _T_1514 & _T_1516; // @[StoreQueue.scala 120:90:@659.4]
  assign _T_1519 = _T_1517 == 1'h0; // @[StoreQueue.scala 120:67:@660.4]
  assign _T_1520 = _T_1444 & _T_1519; // @[StoreQueue.scala 120:64:@661.4]
  assign validEntriesInLoadQ_4 = _T_1437 ? _T_1510 : _T_1520; // @[StoreQueue.scala 119:90:@662.4]
  assign _T_1524 = io_loadHead <= 3'h5; // @[StoreQueue.scala 120:17:@664.4]
  assign _T_1526 = 3'h5 < io_loadTail; // @[StoreQueue.scala 120:35:@665.4]
  assign _T_1527 = _T_1524 & _T_1526; // @[StoreQueue.scala 120:26:@666.4]
  assign _T_1531 = io_loadTail <= 3'h5; // @[StoreQueue.scala 120:81:@668.4]
  assign _T_1533 = 3'h5 < io_loadHead; // @[StoreQueue.scala 120:99:@669.4]
  assign _T_1534 = _T_1531 & _T_1533; // @[StoreQueue.scala 120:90:@670.4]
  assign _T_1536 = _T_1534 == 1'h0; // @[StoreQueue.scala 120:67:@671.4]
  assign _T_1537 = _T_1444 & _T_1536; // @[StoreQueue.scala 120:64:@672.4]
  assign validEntriesInLoadQ_5 = _T_1437 ? _T_1527 : _T_1537; // @[StoreQueue.scala 119:90:@673.4]
  assign _T_1541 = io_loadHead <= 3'h6; // @[StoreQueue.scala 120:17:@675.4]
  assign _T_1543 = 3'h6 < io_loadTail; // @[StoreQueue.scala 120:35:@676.4]
  assign _T_1544 = _T_1541 & _T_1543; // @[StoreQueue.scala 120:26:@677.4]
  assign _T_1548 = io_loadTail <= 3'h6; // @[StoreQueue.scala 120:81:@679.4]
  assign _T_1550 = 3'h6 < io_loadHead; // @[StoreQueue.scala 120:99:@680.4]
  assign _T_1551 = _T_1548 & _T_1550; // @[StoreQueue.scala 120:90:@681.4]
  assign _T_1553 = _T_1551 == 1'h0; // @[StoreQueue.scala 120:67:@682.4]
  assign _T_1554 = _T_1444 & _T_1553; // @[StoreQueue.scala 120:64:@683.4]
  assign validEntriesInLoadQ_6 = _T_1437 ? _T_1544 : _T_1554; // @[StoreQueue.scala 119:90:@684.4]
  assign validEntriesInLoadQ_7 = _T_1437 ? 1'h0 : _T_1444; // @[StoreQueue.scala 119:90:@695.4]
  assign _GEN_241 = 3'h1 == head ? offsetQ_1 : offsetQ_0; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_242 = 3'h2 == head ? offsetQ_2 : _GEN_241; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_243 = 3'h3 == head ? offsetQ_3 : _GEN_242; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_244 = 3'h4 == head ? offsetQ_4 : _GEN_243; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_245 = 3'h5 == head ? offsetQ_5 : _GEN_244; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_246 = 3'h6 == head ? offsetQ_6 : _GEN_245; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_247 = 3'h7 == head ? offsetQ_7 : _GEN_246; // @[StoreQueue.scala 126:96:@705.4]
  assign _T_1589 = io_loadHead <= _GEN_247; // @[StoreQueue.scala 126:96:@705.4]
  assign loadsToCheck_0 = _T_1589 ? _T_1439 : 1'h1; // @[StoreQueue.scala 126:83:@713.4]
  assign _T_1619 = 3'h1 <= _GEN_247; // @[StoreQueue.scala 127:37:@716.4]
  assign _T_1620 = _T_1456 & _T_1619; // @[StoreQueue.scala 127:28:@717.4]
  assign _T_1625 = _GEN_247 < 3'h1; // @[StoreQueue.scala 127:71:@718.4]
  assign _T_1628 = _T_1625 & _T_1465; // @[StoreQueue.scala 127:79:@720.4]
  assign _T_1630 = _T_1628 == 1'h0; // @[StoreQueue.scala 127:55:@721.4]
  assign loadsToCheck_1 = _T_1589 ? _T_1620 : _T_1630; // @[StoreQueue.scala 126:83:@722.4]
  assign _T_1642 = 3'h2 <= _GEN_247; // @[StoreQueue.scala 127:37:@725.4]
  assign _T_1643 = _T_1473 & _T_1642; // @[StoreQueue.scala 127:28:@726.4]
  assign _T_1648 = _GEN_247 < 3'h2; // @[StoreQueue.scala 127:71:@727.4]
  assign _T_1651 = _T_1648 & _T_1482; // @[StoreQueue.scala 127:79:@729.4]
  assign _T_1653 = _T_1651 == 1'h0; // @[StoreQueue.scala 127:55:@730.4]
  assign loadsToCheck_2 = _T_1589 ? _T_1643 : _T_1653; // @[StoreQueue.scala 126:83:@731.4]
  assign _T_1665 = 3'h3 <= _GEN_247; // @[StoreQueue.scala 127:37:@734.4]
  assign _T_1666 = _T_1490 & _T_1665; // @[StoreQueue.scala 127:28:@735.4]
  assign _T_1671 = _GEN_247 < 3'h3; // @[StoreQueue.scala 127:71:@736.4]
  assign _T_1674 = _T_1671 & _T_1499; // @[StoreQueue.scala 127:79:@738.4]
  assign _T_1676 = _T_1674 == 1'h0; // @[StoreQueue.scala 127:55:@739.4]
  assign loadsToCheck_3 = _T_1589 ? _T_1666 : _T_1676; // @[StoreQueue.scala 126:83:@740.4]
  assign _T_1688 = 3'h4 <= _GEN_247; // @[StoreQueue.scala 127:37:@743.4]
  assign _T_1689 = _T_1507 & _T_1688; // @[StoreQueue.scala 127:28:@744.4]
  assign _T_1694 = _GEN_247 < 3'h4; // @[StoreQueue.scala 127:71:@745.4]
  assign _T_1697 = _T_1694 & _T_1516; // @[StoreQueue.scala 127:79:@747.4]
  assign _T_1699 = _T_1697 == 1'h0; // @[StoreQueue.scala 127:55:@748.4]
  assign loadsToCheck_4 = _T_1589 ? _T_1689 : _T_1699; // @[StoreQueue.scala 126:83:@749.4]
  assign _T_1711 = 3'h5 <= _GEN_247; // @[StoreQueue.scala 127:37:@752.4]
  assign _T_1712 = _T_1524 & _T_1711; // @[StoreQueue.scala 127:28:@753.4]
  assign _T_1717 = _GEN_247 < 3'h5; // @[StoreQueue.scala 127:71:@754.4]
  assign _T_1720 = _T_1717 & _T_1533; // @[StoreQueue.scala 127:79:@756.4]
  assign _T_1722 = _T_1720 == 1'h0; // @[StoreQueue.scala 127:55:@757.4]
  assign loadsToCheck_5 = _T_1589 ? _T_1712 : _T_1722; // @[StoreQueue.scala 126:83:@758.4]
  assign _T_1734 = 3'h6 <= _GEN_247; // @[StoreQueue.scala 127:37:@761.4]
  assign _T_1735 = _T_1541 & _T_1734; // @[StoreQueue.scala 127:28:@762.4]
  assign _T_1740 = _GEN_247 < 3'h6; // @[StoreQueue.scala 127:71:@763.4]
  assign _T_1743 = _T_1740 & _T_1550; // @[StoreQueue.scala 127:79:@765.4]
  assign _T_1745 = _T_1743 == 1'h0; // @[StoreQueue.scala 127:55:@766.4]
  assign loadsToCheck_6 = _T_1589 ? _T_1735 : _T_1745; // @[StoreQueue.scala 126:83:@767.4]
  assign _T_1757 = 3'h7 <= _GEN_247; // @[StoreQueue.scala 127:37:@770.4]
  assign loadsToCheck_7 = _T_1589 ? _T_1757 : 1'h1; // @[StoreQueue.scala 126:83:@776.4]
  assign _T_1783 = loadsToCheck_0 & validEntriesInLoadQ_0; // @[StoreQueue.scala 133:16:@786.4]
  assign _GEN_249 = 3'h1 == head ? checkBits_1 : checkBits_0; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_250 = 3'h2 == head ? checkBits_2 : _GEN_249; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_251 = 3'h3 == head ? checkBits_3 : _GEN_250; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_252 = 3'h4 == head ? checkBits_4 : _GEN_251; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_253 = 3'h5 == head ? checkBits_5 : _GEN_252; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_254 = 3'h6 == head ? checkBits_6 : _GEN_253; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_255 = 3'h7 == head ? checkBits_7 : _GEN_254; // @[StoreQueue.scala 133:24:@787.4]
  assign entriesToCheck_0 = _T_1783 & _GEN_255; // @[StoreQueue.scala 133:24:@787.4]
  assign _T_1788 = loadsToCheck_1 & validEntriesInLoadQ_1; // @[StoreQueue.scala 133:16:@788.4]
  assign entriesToCheck_1 = _T_1788 & _GEN_255; // @[StoreQueue.scala 133:24:@789.4]
  assign _T_1793 = loadsToCheck_2 & validEntriesInLoadQ_2; // @[StoreQueue.scala 133:16:@790.4]
  assign entriesToCheck_2 = _T_1793 & _GEN_255; // @[StoreQueue.scala 133:24:@791.4]
  assign _T_1798 = loadsToCheck_3 & validEntriesInLoadQ_3; // @[StoreQueue.scala 133:16:@792.4]
  assign entriesToCheck_3 = _T_1798 & _GEN_255; // @[StoreQueue.scala 133:24:@793.4]
  assign _T_1803 = loadsToCheck_4 & validEntriesInLoadQ_4; // @[StoreQueue.scala 133:16:@794.4]
  assign entriesToCheck_4 = _T_1803 & _GEN_255; // @[StoreQueue.scala 133:24:@795.4]
  assign _T_1808 = loadsToCheck_5 & validEntriesInLoadQ_5; // @[StoreQueue.scala 133:16:@796.4]
  assign entriesToCheck_5 = _T_1808 & _GEN_255; // @[StoreQueue.scala 133:24:@797.4]
  assign _T_1813 = loadsToCheck_6 & validEntriesInLoadQ_6; // @[StoreQueue.scala 133:16:@798.4]
  assign entriesToCheck_6 = _T_1813 & _GEN_255; // @[StoreQueue.scala 133:24:@799.4]
  assign _T_1818 = loadsToCheck_7 & validEntriesInLoadQ_7; // @[StoreQueue.scala 133:16:@800.4]
  assign entriesToCheck_7 = _T_1818 & _GEN_255; // @[StoreQueue.scala 133:24:@801.4]
  assign _T_1850 = entriesToCheck_0 == 1'h0; // @[StoreQueue.scala 140:34:@812.4]
  assign _T_1851 = _T_1850 | io_loadDataDone_0; // @[StoreQueue.scala 140:64:@813.4]
  assign _GEN_257 = 3'h1 == head ? addrQ_1 : addrQ_0; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_258 = 3'h2 == head ? addrQ_2 : _GEN_257; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_259 = 3'h3 == head ? addrQ_3 : _GEN_258; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_260 = 3'h4 == head ? addrQ_4 : _GEN_259; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_261 = 3'h5 == head ? addrQ_5 : _GEN_260; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_262 = 3'h6 == head ? addrQ_6 : _GEN_261; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_263 = 3'h7 == head ? addrQ_7 : _GEN_262; // @[StoreQueue.scala 141:51:@814.4]
  assign _T_1855 = _GEN_263 != io_loadAddressQueue_0; // @[StoreQueue.scala 141:51:@814.4]
  assign _T_1856 = io_loadAddressDone_0 & _T_1855; // @[StoreQueue.scala 141:36:@815.4]
  assign noConflicts_0 = _T_1851 | _T_1856; // @[StoreQueue.scala 140:95:@816.4]
  assign _T_1859 = entriesToCheck_1 == 1'h0; // @[StoreQueue.scala 140:34:@818.4]
  assign _T_1860 = _T_1859 | io_loadDataDone_1; // @[StoreQueue.scala 140:64:@819.4]
  assign _T_1864 = _GEN_263 != io_loadAddressQueue_1; // @[StoreQueue.scala 141:51:@820.4]
  assign _T_1865 = io_loadAddressDone_1 & _T_1864; // @[StoreQueue.scala 141:36:@821.4]
  assign noConflicts_1 = _T_1860 | _T_1865; // @[StoreQueue.scala 140:95:@822.4]
  assign _T_1868 = entriesToCheck_2 == 1'h0; // @[StoreQueue.scala 140:34:@824.4]
  assign _T_1869 = _T_1868 | io_loadDataDone_2; // @[StoreQueue.scala 140:64:@825.4]
  assign _T_1873 = _GEN_263 != io_loadAddressQueue_2; // @[StoreQueue.scala 141:51:@826.4]
  assign _T_1874 = io_loadAddressDone_2 & _T_1873; // @[StoreQueue.scala 141:36:@827.4]
  assign noConflicts_2 = _T_1869 | _T_1874; // @[StoreQueue.scala 140:95:@828.4]
  assign _T_1877 = entriesToCheck_3 == 1'h0; // @[StoreQueue.scala 140:34:@830.4]
  assign _T_1878 = _T_1877 | io_loadDataDone_3; // @[StoreQueue.scala 140:64:@831.4]
  assign _T_1882 = _GEN_263 != io_loadAddressQueue_3; // @[StoreQueue.scala 141:51:@832.4]
  assign _T_1883 = io_loadAddressDone_3 & _T_1882; // @[StoreQueue.scala 141:36:@833.4]
  assign noConflicts_3 = _T_1878 | _T_1883; // @[StoreQueue.scala 140:95:@834.4]
  assign _T_1886 = entriesToCheck_4 == 1'h0; // @[StoreQueue.scala 140:34:@836.4]
  assign _T_1887 = _T_1886 | io_loadDataDone_4; // @[StoreQueue.scala 140:64:@837.4]
  assign _T_1891 = _GEN_263 != io_loadAddressQueue_4; // @[StoreQueue.scala 141:51:@838.4]
  assign _T_1892 = io_loadAddressDone_4 & _T_1891; // @[StoreQueue.scala 141:36:@839.4]
  assign noConflicts_4 = _T_1887 | _T_1892; // @[StoreQueue.scala 140:95:@840.4]
  assign _T_1895 = entriesToCheck_5 == 1'h0; // @[StoreQueue.scala 140:34:@842.4]
  assign _T_1896 = _T_1895 | io_loadDataDone_5; // @[StoreQueue.scala 140:64:@843.4]
  assign _T_1900 = _GEN_263 != io_loadAddressQueue_5; // @[StoreQueue.scala 141:51:@844.4]
  assign _T_1901 = io_loadAddressDone_5 & _T_1900; // @[StoreQueue.scala 141:36:@845.4]
  assign noConflicts_5 = _T_1896 | _T_1901; // @[StoreQueue.scala 140:95:@846.4]
  assign _T_1904 = entriesToCheck_6 == 1'h0; // @[StoreQueue.scala 140:34:@848.4]
  assign _T_1905 = _T_1904 | io_loadDataDone_6; // @[StoreQueue.scala 140:64:@849.4]
  assign _T_1909 = _GEN_263 != io_loadAddressQueue_6; // @[StoreQueue.scala 141:51:@850.4]
  assign _T_1910 = io_loadAddressDone_6 & _T_1909; // @[StoreQueue.scala 141:36:@851.4]
  assign noConflicts_6 = _T_1905 | _T_1910; // @[StoreQueue.scala 140:95:@852.4]
  assign _T_1913 = entriesToCheck_7 == 1'h0; // @[StoreQueue.scala 140:34:@854.4]
  assign _T_1914 = _T_1913 | io_loadDataDone_7; // @[StoreQueue.scala 140:64:@855.4]
  assign _T_1918 = _GEN_263 != io_loadAddressQueue_7; // @[StoreQueue.scala 141:51:@856.4]
  assign _T_1919 = io_loadAddressDone_7 & _T_1918; // @[StoreQueue.scala 141:36:@857.4]
  assign noConflicts_7 = _T_1914 | _T_1919; // @[StoreQueue.scala 140:95:@858.4]
  assign _GEN_265 = 3'h1 == head ? addrKnown_1 : addrKnown_0; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_266 = 3'h2 == head ? addrKnown_2 : _GEN_265; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_267 = 3'h3 == head ? addrKnown_3 : _GEN_266; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_268 = 3'h4 == head ? addrKnown_4 : _GEN_267; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_269 = 3'h5 == head ? addrKnown_5 : _GEN_268; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_270 = 3'h6 == head ? addrKnown_6 : _GEN_269; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_271 = 3'h7 == head ? addrKnown_7 : _GEN_270; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_273 = 3'h1 == head ? dataKnown_1 : dataKnown_0; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_274 = 3'h2 == head ? dataKnown_2 : _GEN_273; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_275 = 3'h3 == head ? dataKnown_3 : _GEN_274; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_276 = 3'h4 == head ? dataKnown_4 : _GEN_275; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_277 = 3'h5 == head ? dataKnown_5 : _GEN_276; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_278 = 3'h6 == head ? dataKnown_6 : _GEN_277; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_279 = 3'h7 == head ? dataKnown_7 : _GEN_278; // @[StoreQueue.scala 154:44:@860.4]
  assign _T_1927 = _GEN_271 & _GEN_279; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_281 = 3'h1 == head ? storeCompleted_1 : storeCompleted_0; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_282 = 3'h2 == head ? storeCompleted_2 : _GEN_281; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_283 = 3'h3 == head ? storeCompleted_3 : _GEN_282; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_284 = 3'h4 == head ? storeCompleted_4 : _GEN_283; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_285 = 3'h5 == head ? storeCompleted_5 : _GEN_284; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_286 = 3'h6 == head ? storeCompleted_6 : _GEN_285; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_287 = 3'h7 == head ? storeCompleted_7 : _GEN_286; // @[StoreQueue.scala 154:66:@861.4]
  assign _T_1932 = _GEN_287 == 1'h0; // @[StoreQueue.scala 154:66:@861.4]
  assign _T_1933 = _T_1927 & _T_1932; // @[StoreQueue.scala 154:63:@862.4]
  assign _T_1936 = noConflicts_0 & noConflicts_1; // @[StoreQueue.scala 154:109:@864.4]
  assign _T_1937 = _T_1936 & noConflicts_2; // @[StoreQueue.scala 154:109:@865.4]
  assign _T_1938 = _T_1937 & noConflicts_3; // @[StoreQueue.scala 154:109:@866.4]
  assign _T_1939 = _T_1938 & noConflicts_4; // @[StoreQueue.scala 154:109:@867.4]
  assign _T_1940 = _T_1939 & noConflicts_5; // @[StoreQueue.scala 154:109:@868.4]
  assign _T_1941 = _T_1940 & noConflicts_6; // @[StoreQueue.scala 154:109:@869.4]
  assign _T_1942 = _T_1941 & noConflicts_7; // @[StoreQueue.scala 154:109:@870.4]
  assign storeRequest = _T_1933 & _T_1942; // @[StoreQueue.scala 154:88:@871.4]
  assign _T_1945 = head == 3'h0; // @[StoreQueue.scala 164:23:@876.6]
  assign _T_1946 = _T_1945 & storeRequest; // @[StoreQueue.scala 164:43:@877.6]
  assign _T_1947 = _T_1946 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@878.6]
  assign _GEN_288 = _T_1947 ? 1'h1 : storeCompleted_0; // @[StoreQueue.scala 164:86:@879.6]
  assign _GEN_289 = initBits_0 ? 1'h0 : _GEN_288; // @[StoreQueue.scala 162:37:@872.4]
  assign _T_1951 = head == 3'h1; // @[StoreQueue.scala 164:23:@886.6]
  assign _T_1952 = _T_1951 & storeRequest; // @[StoreQueue.scala 164:43:@887.6]
  assign _T_1953 = _T_1952 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@888.6]
  assign _GEN_290 = _T_1953 ? 1'h1 : storeCompleted_1; // @[StoreQueue.scala 164:86:@889.6]
  assign _GEN_291 = initBits_1 ? 1'h0 : _GEN_290; // @[StoreQueue.scala 162:37:@882.4]
  assign _T_1957 = head == 3'h2; // @[StoreQueue.scala 164:23:@896.6]
  assign _T_1958 = _T_1957 & storeRequest; // @[StoreQueue.scala 164:43:@897.6]
  assign _T_1959 = _T_1958 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@898.6]
  assign _GEN_292 = _T_1959 ? 1'h1 : storeCompleted_2; // @[StoreQueue.scala 164:86:@899.6]
  assign _GEN_293 = initBits_2 ? 1'h0 : _GEN_292; // @[StoreQueue.scala 162:37:@892.4]
  assign _T_1963 = head == 3'h3; // @[StoreQueue.scala 164:23:@906.6]
  assign _T_1964 = _T_1963 & storeRequest; // @[StoreQueue.scala 164:43:@907.6]
  assign _T_1965 = _T_1964 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@908.6]
  assign _GEN_294 = _T_1965 ? 1'h1 : storeCompleted_3; // @[StoreQueue.scala 164:86:@909.6]
  assign _GEN_295 = initBits_3 ? 1'h0 : _GEN_294; // @[StoreQueue.scala 162:37:@902.4]
  assign _T_1969 = head == 3'h4; // @[StoreQueue.scala 164:23:@916.6]
  assign _T_1970 = _T_1969 & storeRequest; // @[StoreQueue.scala 164:43:@917.6]
  assign _T_1971 = _T_1970 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@918.6]
  assign _GEN_296 = _T_1971 ? 1'h1 : storeCompleted_4; // @[StoreQueue.scala 164:86:@919.6]
  assign _GEN_297 = initBits_4 ? 1'h0 : _GEN_296; // @[StoreQueue.scala 162:37:@912.4]
  assign _T_1975 = head == 3'h5; // @[StoreQueue.scala 164:23:@926.6]
  assign _T_1976 = _T_1975 & storeRequest; // @[StoreQueue.scala 164:43:@927.6]
  assign _T_1977 = _T_1976 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@928.6]
  assign _GEN_298 = _T_1977 ? 1'h1 : storeCompleted_5; // @[StoreQueue.scala 164:86:@929.6]
  assign _GEN_299 = initBits_5 ? 1'h0 : _GEN_298; // @[StoreQueue.scala 162:37:@922.4]
  assign _T_1981 = head == 3'h6; // @[StoreQueue.scala 164:23:@936.6]
  assign _T_1982 = _T_1981 & storeRequest; // @[StoreQueue.scala 164:43:@937.6]
  assign _T_1983 = _T_1982 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@938.6]
  assign _GEN_300 = _T_1983 ? 1'h1 : storeCompleted_6; // @[StoreQueue.scala 164:86:@939.6]
  assign _GEN_301 = initBits_6 ? 1'h0 : _GEN_300; // @[StoreQueue.scala 162:37:@932.4]
  assign _T_1987 = head == 3'h7; // @[StoreQueue.scala 164:23:@946.6]
  assign _T_1988 = _T_1987 & storeRequest; // @[StoreQueue.scala 164:43:@947.6]
  assign _T_1989 = _T_1988 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@948.6]
  assign _GEN_302 = _T_1989 ? 1'h1 : storeCompleted_7; // @[StoreQueue.scala 164:86:@949.6]
  assign _GEN_303 = initBits_7 ? 1'h0 : _GEN_302; // @[StoreQueue.scala 162:37:@942.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[StoreQueue.scala 180:72:@953.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[StoreQueue.scala 180:72:@955.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[StoreQueue.scala 180:72:@957.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[StoreQueue.scala 180:72:@959.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[StoreQueue.scala 180:72:@961.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[StoreQueue.scala 180:72:@963.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[StoreQueue.scala 180:72:@965.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[StoreQueue.scala 180:72:@967.4]
  assign _T_2266 = addrKnown_0 == 1'h0; // @[StoreQueue.scala 192:91:@971.4]
  assign _T_2267 = entriesPorts_0_0 & _T_2266; // @[StoreQueue.scala 192:88:@972.4]
  assign _T_2269 = addrKnown_1 == 1'h0; // @[StoreQueue.scala 192:91:@973.4]
  assign _T_2270 = entriesPorts_0_1 & _T_2269; // @[StoreQueue.scala 192:88:@974.4]
  assign _T_2272 = addrKnown_2 == 1'h0; // @[StoreQueue.scala 192:91:@975.4]
  assign _T_2273 = entriesPorts_0_2 & _T_2272; // @[StoreQueue.scala 192:88:@976.4]
  assign _T_2275 = addrKnown_3 == 1'h0; // @[StoreQueue.scala 192:91:@977.4]
  assign _T_2276 = entriesPorts_0_3 & _T_2275; // @[StoreQueue.scala 192:88:@978.4]
  assign _T_2278 = addrKnown_4 == 1'h0; // @[StoreQueue.scala 192:91:@979.4]
  assign _T_2279 = entriesPorts_0_4 & _T_2278; // @[StoreQueue.scala 192:88:@980.4]
  assign _T_2281 = addrKnown_5 == 1'h0; // @[StoreQueue.scala 192:91:@981.4]
  assign _T_2282 = entriesPorts_0_5 & _T_2281; // @[StoreQueue.scala 192:88:@982.4]
  assign _T_2284 = addrKnown_6 == 1'h0; // @[StoreQueue.scala 192:91:@983.4]
  assign _T_2285 = entriesPorts_0_6 & _T_2284; // @[StoreQueue.scala 192:88:@984.4]
  assign _T_2287 = addrKnown_7 == 1'h0; // @[StoreQueue.scala 192:91:@985.4]
  assign _T_2288 = entriesPorts_0_7 & _T_2287; // @[StoreQueue.scala 192:88:@986.4]
  assign _T_2304 = dataKnown_0 == 1'h0; // @[StoreQueue.scala 193:91:@996.4]
  assign _T_2305 = entriesPorts_0_0 & _T_2304; // @[StoreQueue.scala 193:88:@997.4]
  assign _T_2307 = dataKnown_1 == 1'h0; // @[StoreQueue.scala 193:91:@998.4]
  assign _T_2308 = entriesPorts_0_1 & _T_2307; // @[StoreQueue.scala 193:88:@999.4]
  assign _T_2310 = dataKnown_2 == 1'h0; // @[StoreQueue.scala 193:91:@1000.4]
  assign _T_2311 = entriesPorts_0_2 & _T_2310; // @[StoreQueue.scala 193:88:@1001.4]
  assign _T_2313 = dataKnown_3 == 1'h0; // @[StoreQueue.scala 193:91:@1002.4]
  assign _T_2314 = entriesPorts_0_3 & _T_2313; // @[StoreQueue.scala 193:88:@1003.4]
  assign _T_2316 = dataKnown_4 == 1'h0; // @[StoreQueue.scala 193:91:@1004.4]
  assign _T_2317 = entriesPorts_0_4 & _T_2316; // @[StoreQueue.scala 193:88:@1005.4]
  assign _T_2319 = dataKnown_5 == 1'h0; // @[StoreQueue.scala 193:91:@1006.4]
  assign _T_2320 = entriesPorts_0_5 & _T_2319; // @[StoreQueue.scala 193:88:@1007.4]
  assign _T_2322 = dataKnown_6 == 1'h0; // @[StoreQueue.scala 193:91:@1008.4]
  assign _T_2323 = entriesPorts_0_6 & _T_2322; // @[StoreQueue.scala 193:88:@1009.4]
  assign _T_2325 = dataKnown_7 == 1'h0; // @[StoreQueue.scala 193:91:@1010.4]
  assign _T_2326 = entriesPorts_0_7 & _T_2325; // @[StoreQueue.scala 193:88:@1011.4]
  assign _T_2343 = 8'h1 << head; // @[OneHot.scala 52:12:@1022.4]
  assign _T_2345 = _T_2343[0]; // @[util.scala 33:60:@1024.4]
  assign _T_2346 = _T_2343[1]; // @[util.scala 33:60:@1025.4]
  assign _T_2347 = _T_2343[2]; // @[util.scala 33:60:@1026.4]
  assign _T_2348 = _T_2343[3]; // @[util.scala 33:60:@1027.4]
  assign _T_2349 = _T_2343[4]; // @[util.scala 33:60:@1028.4]
  assign _T_2350 = _T_2343[5]; // @[util.scala 33:60:@1029.4]
  assign _T_2351 = _T_2343[6]; // @[util.scala 33:60:@1030.4]
  assign _T_2352 = _T_2343[7]; // @[util.scala 33:60:@1031.4]
  assign _T_2377 = _T_2288 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1041.4]
  assign _T_2378 = _T_2285 ? 8'h40 : _T_2377; // @[Mux.scala 31:69:@1042.4]
  assign _T_2379 = _T_2282 ? 8'h20 : _T_2378; // @[Mux.scala 31:69:@1043.4]
  assign _T_2380 = _T_2279 ? 8'h10 : _T_2379; // @[Mux.scala 31:69:@1044.4]
  assign _T_2381 = _T_2276 ? 8'h8 : _T_2380; // @[Mux.scala 31:69:@1045.4]
  assign _T_2382 = _T_2273 ? 8'h4 : _T_2381; // @[Mux.scala 31:69:@1046.4]
  assign _T_2383 = _T_2270 ? 8'h2 : _T_2382; // @[Mux.scala 31:69:@1047.4]
  assign _T_2384 = _T_2267 ? 8'h1 : _T_2383; // @[Mux.scala 31:69:@1048.4]
  assign _T_2385 = _T_2384[0]; // @[OneHot.scala 66:30:@1049.4]
  assign _T_2386 = _T_2384[1]; // @[OneHot.scala 66:30:@1050.4]
  assign _T_2387 = _T_2384[2]; // @[OneHot.scala 66:30:@1051.4]
  assign _T_2388 = _T_2384[3]; // @[OneHot.scala 66:30:@1052.4]
  assign _T_2389 = _T_2384[4]; // @[OneHot.scala 66:30:@1053.4]
  assign _T_2390 = _T_2384[5]; // @[OneHot.scala 66:30:@1054.4]
  assign _T_2391 = _T_2384[6]; // @[OneHot.scala 66:30:@1055.4]
  assign _T_2392 = _T_2384[7]; // @[OneHot.scala 66:30:@1056.4]
  assign _T_2417 = _T_2267 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1066.4]
  assign _T_2418 = _T_2288 ? 8'h40 : _T_2417; // @[Mux.scala 31:69:@1067.4]
  assign _T_2419 = _T_2285 ? 8'h20 : _T_2418; // @[Mux.scala 31:69:@1068.4]
  assign _T_2420 = _T_2282 ? 8'h10 : _T_2419; // @[Mux.scala 31:69:@1069.4]
  assign _T_2421 = _T_2279 ? 8'h8 : _T_2420; // @[Mux.scala 31:69:@1070.4]
  assign _T_2422 = _T_2276 ? 8'h4 : _T_2421; // @[Mux.scala 31:69:@1071.4]
  assign _T_2423 = _T_2273 ? 8'h2 : _T_2422; // @[Mux.scala 31:69:@1072.4]
  assign _T_2424 = _T_2270 ? 8'h1 : _T_2423; // @[Mux.scala 31:69:@1073.4]
  assign _T_2425 = _T_2424[0]; // @[OneHot.scala 66:30:@1074.4]
  assign _T_2426 = _T_2424[1]; // @[OneHot.scala 66:30:@1075.4]
  assign _T_2427 = _T_2424[2]; // @[OneHot.scala 66:30:@1076.4]
  assign _T_2428 = _T_2424[3]; // @[OneHot.scala 66:30:@1077.4]
  assign _T_2429 = _T_2424[4]; // @[OneHot.scala 66:30:@1078.4]
  assign _T_2430 = _T_2424[5]; // @[OneHot.scala 66:30:@1079.4]
  assign _T_2431 = _T_2424[6]; // @[OneHot.scala 66:30:@1080.4]
  assign _T_2432 = _T_2424[7]; // @[OneHot.scala 66:30:@1081.4]
  assign _T_2457 = _T_2270 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1091.4]
  assign _T_2458 = _T_2267 ? 8'h40 : _T_2457; // @[Mux.scala 31:69:@1092.4]
  assign _T_2459 = _T_2288 ? 8'h20 : _T_2458; // @[Mux.scala 31:69:@1093.4]
  assign _T_2460 = _T_2285 ? 8'h10 : _T_2459; // @[Mux.scala 31:69:@1094.4]
  assign _T_2461 = _T_2282 ? 8'h8 : _T_2460; // @[Mux.scala 31:69:@1095.4]
  assign _T_2462 = _T_2279 ? 8'h4 : _T_2461; // @[Mux.scala 31:69:@1096.4]
  assign _T_2463 = _T_2276 ? 8'h2 : _T_2462; // @[Mux.scala 31:69:@1097.4]
  assign _T_2464 = _T_2273 ? 8'h1 : _T_2463; // @[Mux.scala 31:69:@1098.4]
  assign _T_2465 = _T_2464[0]; // @[OneHot.scala 66:30:@1099.4]
  assign _T_2466 = _T_2464[1]; // @[OneHot.scala 66:30:@1100.4]
  assign _T_2467 = _T_2464[2]; // @[OneHot.scala 66:30:@1101.4]
  assign _T_2468 = _T_2464[3]; // @[OneHot.scala 66:30:@1102.4]
  assign _T_2469 = _T_2464[4]; // @[OneHot.scala 66:30:@1103.4]
  assign _T_2470 = _T_2464[5]; // @[OneHot.scala 66:30:@1104.4]
  assign _T_2471 = _T_2464[6]; // @[OneHot.scala 66:30:@1105.4]
  assign _T_2472 = _T_2464[7]; // @[OneHot.scala 66:30:@1106.4]
  assign _T_2497 = _T_2273 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1116.4]
  assign _T_2498 = _T_2270 ? 8'h40 : _T_2497; // @[Mux.scala 31:69:@1117.4]
  assign _T_2499 = _T_2267 ? 8'h20 : _T_2498; // @[Mux.scala 31:69:@1118.4]
  assign _T_2500 = _T_2288 ? 8'h10 : _T_2499; // @[Mux.scala 31:69:@1119.4]
  assign _T_2501 = _T_2285 ? 8'h8 : _T_2500; // @[Mux.scala 31:69:@1120.4]
  assign _T_2502 = _T_2282 ? 8'h4 : _T_2501; // @[Mux.scala 31:69:@1121.4]
  assign _T_2503 = _T_2279 ? 8'h2 : _T_2502; // @[Mux.scala 31:69:@1122.4]
  assign _T_2504 = _T_2276 ? 8'h1 : _T_2503; // @[Mux.scala 31:69:@1123.4]
  assign _T_2505 = _T_2504[0]; // @[OneHot.scala 66:30:@1124.4]
  assign _T_2506 = _T_2504[1]; // @[OneHot.scala 66:30:@1125.4]
  assign _T_2507 = _T_2504[2]; // @[OneHot.scala 66:30:@1126.4]
  assign _T_2508 = _T_2504[3]; // @[OneHot.scala 66:30:@1127.4]
  assign _T_2509 = _T_2504[4]; // @[OneHot.scala 66:30:@1128.4]
  assign _T_2510 = _T_2504[5]; // @[OneHot.scala 66:30:@1129.4]
  assign _T_2511 = _T_2504[6]; // @[OneHot.scala 66:30:@1130.4]
  assign _T_2512 = _T_2504[7]; // @[OneHot.scala 66:30:@1131.4]
  assign _T_2537 = _T_2276 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1141.4]
  assign _T_2538 = _T_2273 ? 8'h40 : _T_2537; // @[Mux.scala 31:69:@1142.4]
  assign _T_2539 = _T_2270 ? 8'h20 : _T_2538; // @[Mux.scala 31:69:@1143.4]
  assign _T_2540 = _T_2267 ? 8'h10 : _T_2539; // @[Mux.scala 31:69:@1144.4]
  assign _T_2541 = _T_2288 ? 8'h8 : _T_2540; // @[Mux.scala 31:69:@1145.4]
  assign _T_2542 = _T_2285 ? 8'h4 : _T_2541; // @[Mux.scala 31:69:@1146.4]
  assign _T_2543 = _T_2282 ? 8'h2 : _T_2542; // @[Mux.scala 31:69:@1147.4]
  assign _T_2544 = _T_2279 ? 8'h1 : _T_2543; // @[Mux.scala 31:69:@1148.4]
  assign _T_2545 = _T_2544[0]; // @[OneHot.scala 66:30:@1149.4]
  assign _T_2546 = _T_2544[1]; // @[OneHot.scala 66:30:@1150.4]
  assign _T_2547 = _T_2544[2]; // @[OneHot.scala 66:30:@1151.4]
  assign _T_2548 = _T_2544[3]; // @[OneHot.scala 66:30:@1152.4]
  assign _T_2549 = _T_2544[4]; // @[OneHot.scala 66:30:@1153.4]
  assign _T_2550 = _T_2544[5]; // @[OneHot.scala 66:30:@1154.4]
  assign _T_2551 = _T_2544[6]; // @[OneHot.scala 66:30:@1155.4]
  assign _T_2552 = _T_2544[7]; // @[OneHot.scala 66:30:@1156.4]
  assign _T_2577 = _T_2279 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1166.4]
  assign _T_2578 = _T_2276 ? 8'h40 : _T_2577; // @[Mux.scala 31:69:@1167.4]
  assign _T_2579 = _T_2273 ? 8'h20 : _T_2578; // @[Mux.scala 31:69:@1168.4]
  assign _T_2580 = _T_2270 ? 8'h10 : _T_2579; // @[Mux.scala 31:69:@1169.4]
  assign _T_2581 = _T_2267 ? 8'h8 : _T_2580; // @[Mux.scala 31:69:@1170.4]
  assign _T_2582 = _T_2288 ? 8'h4 : _T_2581; // @[Mux.scala 31:69:@1171.4]
  assign _T_2583 = _T_2285 ? 8'h2 : _T_2582; // @[Mux.scala 31:69:@1172.4]
  assign _T_2584 = _T_2282 ? 8'h1 : _T_2583; // @[Mux.scala 31:69:@1173.4]
  assign _T_2585 = _T_2584[0]; // @[OneHot.scala 66:30:@1174.4]
  assign _T_2586 = _T_2584[1]; // @[OneHot.scala 66:30:@1175.4]
  assign _T_2587 = _T_2584[2]; // @[OneHot.scala 66:30:@1176.4]
  assign _T_2588 = _T_2584[3]; // @[OneHot.scala 66:30:@1177.4]
  assign _T_2589 = _T_2584[4]; // @[OneHot.scala 66:30:@1178.4]
  assign _T_2590 = _T_2584[5]; // @[OneHot.scala 66:30:@1179.4]
  assign _T_2591 = _T_2584[6]; // @[OneHot.scala 66:30:@1180.4]
  assign _T_2592 = _T_2584[7]; // @[OneHot.scala 66:30:@1181.4]
  assign _T_2617 = _T_2282 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1191.4]
  assign _T_2618 = _T_2279 ? 8'h40 : _T_2617; // @[Mux.scala 31:69:@1192.4]
  assign _T_2619 = _T_2276 ? 8'h20 : _T_2618; // @[Mux.scala 31:69:@1193.4]
  assign _T_2620 = _T_2273 ? 8'h10 : _T_2619; // @[Mux.scala 31:69:@1194.4]
  assign _T_2621 = _T_2270 ? 8'h8 : _T_2620; // @[Mux.scala 31:69:@1195.4]
  assign _T_2622 = _T_2267 ? 8'h4 : _T_2621; // @[Mux.scala 31:69:@1196.4]
  assign _T_2623 = _T_2288 ? 8'h2 : _T_2622; // @[Mux.scala 31:69:@1197.4]
  assign _T_2624 = _T_2285 ? 8'h1 : _T_2623; // @[Mux.scala 31:69:@1198.4]
  assign _T_2625 = _T_2624[0]; // @[OneHot.scala 66:30:@1199.4]
  assign _T_2626 = _T_2624[1]; // @[OneHot.scala 66:30:@1200.4]
  assign _T_2627 = _T_2624[2]; // @[OneHot.scala 66:30:@1201.4]
  assign _T_2628 = _T_2624[3]; // @[OneHot.scala 66:30:@1202.4]
  assign _T_2629 = _T_2624[4]; // @[OneHot.scala 66:30:@1203.4]
  assign _T_2630 = _T_2624[5]; // @[OneHot.scala 66:30:@1204.4]
  assign _T_2631 = _T_2624[6]; // @[OneHot.scala 66:30:@1205.4]
  assign _T_2632 = _T_2624[7]; // @[OneHot.scala 66:30:@1206.4]
  assign _T_2657 = _T_2285 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1216.4]
  assign _T_2658 = _T_2282 ? 8'h40 : _T_2657; // @[Mux.scala 31:69:@1217.4]
  assign _T_2659 = _T_2279 ? 8'h20 : _T_2658; // @[Mux.scala 31:69:@1218.4]
  assign _T_2660 = _T_2276 ? 8'h10 : _T_2659; // @[Mux.scala 31:69:@1219.4]
  assign _T_2661 = _T_2273 ? 8'h8 : _T_2660; // @[Mux.scala 31:69:@1220.4]
  assign _T_2662 = _T_2270 ? 8'h4 : _T_2661; // @[Mux.scala 31:69:@1221.4]
  assign _T_2663 = _T_2267 ? 8'h2 : _T_2662; // @[Mux.scala 31:69:@1222.4]
  assign _T_2664 = _T_2288 ? 8'h1 : _T_2663; // @[Mux.scala 31:69:@1223.4]
  assign _T_2665 = _T_2664[0]; // @[OneHot.scala 66:30:@1224.4]
  assign _T_2666 = _T_2664[1]; // @[OneHot.scala 66:30:@1225.4]
  assign _T_2667 = _T_2664[2]; // @[OneHot.scala 66:30:@1226.4]
  assign _T_2668 = _T_2664[3]; // @[OneHot.scala 66:30:@1227.4]
  assign _T_2669 = _T_2664[4]; // @[OneHot.scala 66:30:@1228.4]
  assign _T_2670 = _T_2664[5]; // @[OneHot.scala 66:30:@1229.4]
  assign _T_2671 = _T_2664[6]; // @[OneHot.scala 66:30:@1230.4]
  assign _T_2672 = _T_2664[7]; // @[OneHot.scala 66:30:@1231.4]
  assign _T_2713 = {_T_2392,_T_2391,_T_2390,_T_2389,_T_2388,_T_2387,_T_2386,_T_2385}; // @[Mux.scala 19:72:@1247.4]
  assign _T_2715 = _T_2345 ? _T_2713 : 8'h0; // @[Mux.scala 19:72:@1248.4]
  assign _T_2722 = {_T_2431,_T_2430,_T_2429,_T_2428,_T_2427,_T_2426,_T_2425,_T_2432}; // @[Mux.scala 19:72:@1255.4]
  assign _T_2724 = _T_2346 ? _T_2722 : 8'h0; // @[Mux.scala 19:72:@1256.4]
  assign _T_2731 = {_T_2470,_T_2469,_T_2468,_T_2467,_T_2466,_T_2465,_T_2472,_T_2471}; // @[Mux.scala 19:72:@1263.4]
  assign _T_2733 = _T_2347 ? _T_2731 : 8'h0; // @[Mux.scala 19:72:@1264.4]
  assign _T_2740 = {_T_2509,_T_2508,_T_2507,_T_2506,_T_2505,_T_2512,_T_2511,_T_2510}; // @[Mux.scala 19:72:@1271.4]
  assign _T_2742 = _T_2348 ? _T_2740 : 8'h0; // @[Mux.scala 19:72:@1272.4]
  assign _T_2749 = {_T_2548,_T_2547,_T_2546,_T_2545,_T_2552,_T_2551,_T_2550,_T_2549}; // @[Mux.scala 19:72:@1279.4]
  assign _T_2751 = _T_2349 ? _T_2749 : 8'h0; // @[Mux.scala 19:72:@1280.4]
  assign _T_2758 = {_T_2587,_T_2586,_T_2585,_T_2592,_T_2591,_T_2590,_T_2589,_T_2588}; // @[Mux.scala 19:72:@1287.4]
  assign _T_2760 = _T_2350 ? _T_2758 : 8'h0; // @[Mux.scala 19:72:@1288.4]
  assign _T_2767 = {_T_2626,_T_2625,_T_2632,_T_2631,_T_2630,_T_2629,_T_2628,_T_2627}; // @[Mux.scala 19:72:@1295.4]
  assign _T_2769 = _T_2351 ? _T_2767 : 8'h0; // @[Mux.scala 19:72:@1296.4]
  assign _T_2776 = {_T_2665,_T_2672,_T_2671,_T_2670,_T_2669,_T_2668,_T_2667,_T_2666}; // @[Mux.scala 19:72:@1303.4]
  assign _T_2778 = _T_2352 ? _T_2776 : 8'h0; // @[Mux.scala 19:72:@1304.4]
  assign _T_2779 = _T_2715 | _T_2724; // @[Mux.scala 19:72:@1305.4]
  assign _T_2780 = _T_2779 | _T_2733; // @[Mux.scala 19:72:@1306.4]
  assign _T_2781 = _T_2780 | _T_2742; // @[Mux.scala 19:72:@1307.4]
  assign _T_2782 = _T_2781 | _T_2751; // @[Mux.scala 19:72:@1308.4]
  assign _T_2783 = _T_2782 | _T_2760; // @[Mux.scala 19:72:@1309.4]
  assign _T_2784 = _T_2783 | _T_2769; // @[Mux.scala 19:72:@1310.4]
  assign _T_2785 = _T_2784 | _T_2778; // @[Mux.scala 19:72:@1311.4]
  assign inputAddrPriorityPorts_0_0 = _T_2785[0]; // @[Mux.scala 19:72:@1315.4]
  assign inputAddrPriorityPorts_0_1 = _T_2785[1]; // @[Mux.scala 19:72:@1317.4]
  assign inputAddrPriorityPorts_0_2 = _T_2785[2]; // @[Mux.scala 19:72:@1319.4]
  assign inputAddrPriorityPorts_0_3 = _T_2785[3]; // @[Mux.scala 19:72:@1321.4]
  assign inputAddrPriorityPorts_0_4 = _T_2785[4]; // @[Mux.scala 19:72:@1323.4]
  assign inputAddrPriorityPorts_0_5 = _T_2785[5]; // @[Mux.scala 19:72:@1325.4]
  assign inputAddrPriorityPorts_0_6 = _T_2785[6]; // @[Mux.scala 19:72:@1327.4]
  assign inputAddrPriorityPorts_0_7 = _T_2785[7]; // @[Mux.scala 19:72:@1329.4]
  assign _T_2899 = _T_2326 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1359.4]
  assign _T_2900 = _T_2323 ? 8'h40 : _T_2899; // @[Mux.scala 31:69:@1360.4]
  assign _T_2901 = _T_2320 ? 8'h20 : _T_2900; // @[Mux.scala 31:69:@1361.4]
  assign _T_2902 = _T_2317 ? 8'h10 : _T_2901; // @[Mux.scala 31:69:@1362.4]
  assign _T_2903 = _T_2314 ? 8'h8 : _T_2902; // @[Mux.scala 31:69:@1363.4]
  assign _T_2904 = _T_2311 ? 8'h4 : _T_2903; // @[Mux.scala 31:69:@1364.4]
  assign _T_2905 = _T_2308 ? 8'h2 : _T_2904; // @[Mux.scala 31:69:@1365.4]
  assign _T_2906 = _T_2305 ? 8'h1 : _T_2905; // @[Mux.scala 31:69:@1366.4]
  assign _T_2907 = _T_2906[0]; // @[OneHot.scala 66:30:@1367.4]
  assign _T_2908 = _T_2906[1]; // @[OneHot.scala 66:30:@1368.4]
  assign _T_2909 = _T_2906[2]; // @[OneHot.scala 66:30:@1369.4]
  assign _T_2910 = _T_2906[3]; // @[OneHot.scala 66:30:@1370.4]
  assign _T_2911 = _T_2906[4]; // @[OneHot.scala 66:30:@1371.4]
  assign _T_2912 = _T_2906[5]; // @[OneHot.scala 66:30:@1372.4]
  assign _T_2913 = _T_2906[6]; // @[OneHot.scala 66:30:@1373.4]
  assign _T_2914 = _T_2906[7]; // @[OneHot.scala 66:30:@1374.4]
  assign _T_2939 = _T_2305 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1384.4]
  assign _T_2940 = _T_2326 ? 8'h40 : _T_2939; // @[Mux.scala 31:69:@1385.4]
  assign _T_2941 = _T_2323 ? 8'h20 : _T_2940; // @[Mux.scala 31:69:@1386.4]
  assign _T_2942 = _T_2320 ? 8'h10 : _T_2941; // @[Mux.scala 31:69:@1387.4]
  assign _T_2943 = _T_2317 ? 8'h8 : _T_2942; // @[Mux.scala 31:69:@1388.4]
  assign _T_2944 = _T_2314 ? 8'h4 : _T_2943; // @[Mux.scala 31:69:@1389.4]
  assign _T_2945 = _T_2311 ? 8'h2 : _T_2944; // @[Mux.scala 31:69:@1390.4]
  assign _T_2946 = _T_2308 ? 8'h1 : _T_2945; // @[Mux.scala 31:69:@1391.4]
  assign _T_2947 = _T_2946[0]; // @[OneHot.scala 66:30:@1392.4]
  assign _T_2948 = _T_2946[1]; // @[OneHot.scala 66:30:@1393.4]
  assign _T_2949 = _T_2946[2]; // @[OneHot.scala 66:30:@1394.4]
  assign _T_2950 = _T_2946[3]; // @[OneHot.scala 66:30:@1395.4]
  assign _T_2951 = _T_2946[4]; // @[OneHot.scala 66:30:@1396.4]
  assign _T_2952 = _T_2946[5]; // @[OneHot.scala 66:30:@1397.4]
  assign _T_2953 = _T_2946[6]; // @[OneHot.scala 66:30:@1398.4]
  assign _T_2954 = _T_2946[7]; // @[OneHot.scala 66:30:@1399.4]
  assign _T_2979 = _T_2308 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1409.4]
  assign _T_2980 = _T_2305 ? 8'h40 : _T_2979; // @[Mux.scala 31:69:@1410.4]
  assign _T_2981 = _T_2326 ? 8'h20 : _T_2980; // @[Mux.scala 31:69:@1411.4]
  assign _T_2982 = _T_2323 ? 8'h10 : _T_2981; // @[Mux.scala 31:69:@1412.4]
  assign _T_2983 = _T_2320 ? 8'h8 : _T_2982; // @[Mux.scala 31:69:@1413.4]
  assign _T_2984 = _T_2317 ? 8'h4 : _T_2983; // @[Mux.scala 31:69:@1414.4]
  assign _T_2985 = _T_2314 ? 8'h2 : _T_2984; // @[Mux.scala 31:69:@1415.4]
  assign _T_2986 = _T_2311 ? 8'h1 : _T_2985; // @[Mux.scala 31:69:@1416.4]
  assign _T_2987 = _T_2986[0]; // @[OneHot.scala 66:30:@1417.4]
  assign _T_2988 = _T_2986[1]; // @[OneHot.scala 66:30:@1418.4]
  assign _T_2989 = _T_2986[2]; // @[OneHot.scala 66:30:@1419.4]
  assign _T_2990 = _T_2986[3]; // @[OneHot.scala 66:30:@1420.4]
  assign _T_2991 = _T_2986[4]; // @[OneHot.scala 66:30:@1421.4]
  assign _T_2992 = _T_2986[5]; // @[OneHot.scala 66:30:@1422.4]
  assign _T_2993 = _T_2986[6]; // @[OneHot.scala 66:30:@1423.4]
  assign _T_2994 = _T_2986[7]; // @[OneHot.scala 66:30:@1424.4]
  assign _T_3019 = _T_2311 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1434.4]
  assign _T_3020 = _T_2308 ? 8'h40 : _T_3019; // @[Mux.scala 31:69:@1435.4]
  assign _T_3021 = _T_2305 ? 8'h20 : _T_3020; // @[Mux.scala 31:69:@1436.4]
  assign _T_3022 = _T_2326 ? 8'h10 : _T_3021; // @[Mux.scala 31:69:@1437.4]
  assign _T_3023 = _T_2323 ? 8'h8 : _T_3022; // @[Mux.scala 31:69:@1438.4]
  assign _T_3024 = _T_2320 ? 8'h4 : _T_3023; // @[Mux.scala 31:69:@1439.4]
  assign _T_3025 = _T_2317 ? 8'h2 : _T_3024; // @[Mux.scala 31:69:@1440.4]
  assign _T_3026 = _T_2314 ? 8'h1 : _T_3025; // @[Mux.scala 31:69:@1441.4]
  assign _T_3027 = _T_3026[0]; // @[OneHot.scala 66:30:@1442.4]
  assign _T_3028 = _T_3026[1]; // @[OneHot.scala 66:30:@1443.4]
  assign _T_3029 = _T_3026[2]; // @[OneHot.scala 66:30:@1444.4]
  assign _T_3030 = _T_3026[3]; // @[OneHot.scala 66:30:@1445.4]
  assign _T_3031 = _T_3026[4]; // @[OneHot.scala 66:30:@1446.4]
  assign _T_3032 = _T_3026[5]; // @[OneHot.scala 66:30:@1447.4]
  assign _T_3033 = _T_3026[6]; // @[OneHot.scala 66:30:@1448.4]
  assign _T_3034 = _T_3026[7]; // @[OneHot.scala 66:30:@1449.4]
  assign _T_3059 = _T_2314 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1459.4]
  assign _T_3060 = _T_2311 ? 8'h40 : _T_3059; // @[Mux.scala 31:69:@1460.4]
  assign _T_3061 = _T_2308 ? 8'h20 : _T_3060; // @[Mux.scala 31:69:@1461.4]
  assign _T_3062 = _T_2305 ? 8'h10 : _T_3061; // @[Mux.scala 31:69:@1462.4]
  assign _T_3063 = _T_2326 ? 8'h8 : _T_3062; // @[Mux.scala 31:69:@1463.4]
  assign _T_3064 = _T_2323 ? 8'h4 : _T_3063; // @[Mux.scala 31:69:@1464.4]
  assign _T_3065 = _T_2320 ? 8'h2 : _T_3064; // @[Mux.scala 31:69:@1465.4]
  assign _T_3066 = _T_2317 ? 8'h1 : _T_3065; // @[Mux.scala 31:69:@1466.4]
  assign _T_3067 = _T_3066[0]; // @[OneHot.scala 66:30:@1467.4]
  assign _T_3068 = _T_3066[1]; // @[OneHot.scala 66:30:@1468.4]
  assign _T_3069 = _T_3066[2]; // @[OneHot.scala 66:30:@1469.4]
  assign _T_3070 = _T_3066[3]; // @[OneHot.scala 66:30:@1470.4]
  assign _T_3071 = _T_3066[4]; // @[OneHot.scala 66:30:@1471.4]
  assign _T_3072 = _T_3066[5]; // @[OneHot.scala 66:30:@1472.4]
  assign _T_3073 = _T_3066[6]; // @[OneHot.scala 66:30:@1473.4]
  assign _T_3074 = _T_3066[7]; // @[OneHot.scala 66:30:@1474.4]
  assign _T_3099 = _T_2317 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1484.4]
  assign _T_3100 = _T_2314 ? 8'h40 : _T_3099; // @[Mux.scala 31:69:@1485.4]
  assign _T_3101 = _T_2311 ? 8'h20 : _T_3100; // @[Mux.scala 31:69:@1486.4]
  assign _T_3102 = _T_2308 ? 8'h10 : _T_3101; // @[Mux.scala 31:69:@1487.4]
  assign _T_3103 = _T_2305 ? 8'h8 : _T_3102; // @[Mux.scala 31:69:@1488.4]
  assign _T_3104 = _T_2326 ? 8'h4 : _T_3103; // @[Mux.scala 31:69:@1489.4]
  assign _T_3105 = _T_2323 ? 8'h2 : _T_3104; // @[Mux.scala 31:69:@1490.4]
  assign _T_3106 = _T_2320 ? 8'h1 : _T_3105; // @[Mux.scala 31:69:@1491.4]
  assign _T_3107 = _T_3106[0]; // @[OneHot.scala 66:30:@1492.4]
  assign _T_3108 = _T_3106[1]; // @[OneHot.scala 66:30:@1493.4]
  assign _T_3109 = _T_3106[2]; // @[OneHot.scala 66:30:@1494.4]
  assign _T_3110 = _T_3106[3]; // @[OneHot.scala 66:30:@1495.4]
  assign _T_3111 = _T_3106[4]; // @[OneHot.scala 66:30:@1496.4]
  assign _T_3112 = _T_3106[5]; // @[OneHot.scala 66:30:@1497.4]
  assign _T_3113 = _T_3106[6]; // @[OneHot.scala 66:30:@1498.4]
  assign _T_3114 = _T_3106[7]; // @[OneHot.scala 66:30:@1499.4]
  assign _T_3139 = _T_2320 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1509.4]
  assign _T_3140 = _T_2317 ? 8'h40 : _T_3139; // @[Mux.scala 31:69:@1510.4]
  assign _T_3141 = _T_2314 ? 8'h20 : _T_3140; // @[Mux.scala 31:69:@1511.4]
  assign _T_3142 = _T_2311 ? 8'h10 : _T_3141; // @[Mux.scala 31:69:@1512.4]
  assign _T_3143 = _T_2308 ? 8'h8 : _T_3142; // @[Mux.scala 31:69:@1513.4]
  assign _T_3144 = _T_2305 ? 8'h4 : _T_3143; // @[Mux.scala 31:69:@1514.4]
  assign _T_3145 = _T_2326 ? 8'h2 : _T_3144; // @[Mux.scala 31:69:@1515.4]
  assign _T_3146 = _T_2323 ? 8'h1 : _T_3145; // @[Mux.scala 31:69:@1516.4]
  assign _T_3147 = _T_3146[0]; // @[OneHot.scala 66:30:@1517.4]
  assign _T_3148 = _T_3146[1]; // @[OneHot.scala 66:30:@1518.4]
  assign _T_3149 = _T_3146[2]; // @[OneHot.scala 66:30:@1519.4]
  assign _T_3150 = _T_3146[3]; // @[OneHot.scala 66:30:@1520.4]
  assign _T_3151 = _T_3146[4]; // @[OneHot.scala 66:30:@1521.4]
  assign _T_3152 = _T_3146[5]; // @[OneHot.scala 66:30:@1522.4]
  assign _T_3153 = _T_3146[6]; // @[OneHot.scala 66:30:@1523.4]
  assign _T_3154 = _T_3146[7]; // @[OneHot.scala 66:30:@1524.4]
  assign _T_3179 = _T_2323 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1534.4]
  assign _T_3180 = _T_2320 ? 8'h40 : _T_3179; // @[Mux.scala 31:69:@1535.4]
  assign _T_3181 = _T_2317 ? 8'h20 : _T_3180; // @[Mux.scala 31:69:@1536.4]
  assign _T_3182 = _T_2314 ? 8'h10 : _T_3181; // @[Mux.scala 31:69:@1537.4]
  assign _T_3183 = _T_2311 ? 8'h8 : _T_3182; // @[Mux.scala 31:69:@1538.4]
  assign _T_3184 = _T_2308 ? 8'h4 : _T_3183; // @[Mux.scala 31:69:@1539.4]
  assign _T_3185 = _T_2305 ? 8'h2 : _T_3184; // @[Mux.scala 31:69:@1540.4]
  assign _T_3186 = _T_2326 ? 8'h1 : _T_3185; // @[Mux.scala 31:69:@1541.4]
  assign _T_3187 = _T_3186[0]; // @[OneHot.scala 66:30:@1542.4]
  assign _T_3188 = _T_3186[1]; // @[OneHot.scala 66:30:@1543.4]
  assign _T_3189 = _T_3186[2]; // @[OneHot.scala 66:30:@1544.4]
  assign _T_3190 = _T_3186[3]; // @[OneHot.scala 66:30:@1545.4]
  assign _T_3191 = _T_3186[4]; // @[OneHot.scala 66:30:@1546.4]
  assign _T_3192 = _T_3186[5]; // @[OneHot.scala 66:30:@1547.4]
  assign _T_3193 = _T_3186[6]; // @[OneHot.scala 66:30:@1548.4]
  assign _T_3194 = _T_3186[7]; // @[OneHot.scala 66:30:@1549.4]
  assign _T_3235 = {_T_2914,_T_2913,_T_2912,_T_2911,_T_2910,_T_2909,_T_2908,_T_2907}; // @[Mux.scala 19:72:@1565.4]
  assign _T_3237 = _T_2345 ? _T_3235 : 8'h0; // @[Mux.scala 19:72:@1566.4]
  assign _T_3244 = {_T_2953,_T_2952,_T_2951,_T_2950,_T_2949,_T_2948,_T_2947,_T_2954}; // @[Mux.scala 19:72:@1573.4]
  assign _T_3246 = _T_2346 ? _T_3244 : 8'h0; // @[Mux.scala 19:72:@1574.4]
  assign _T_3253 = {_T_2992,_T_2991,_T_2990,_T_2989,_T_2988,_T_2987,_T_2994,_T_2993}; // @[Mux.scala 19:72:@1581.4]
  assign _T_3255 = _T_2347 ? _T_3253 : 8'h0; // @[Mux.scala 19:72:@1582.4]
  assign _T_3262 = {_T_3031,_T_3030,_T_3029,_T_3028,_T_3027,_T_3034,_T_3033,_T_3032}; // @[Mux.scala 19:72:@1589.4]
  assign _T_3264 = _T_2348 ? _T_3262 : 8'h0; // @[Mux.scala 19:72:@1590.4]
  assign _T_3271 = {_T_3070,_T_3069,_T_3068,_T_3067,_T_3074,_T_3073,_T_3072,_T_3071}; // @[Mux.scala 19:72:@1597.4]
  assign _T_3273 = _T_2349 ? _T_3271 : 8'h0; // @[Mux.scala 19:72:@1598.4]
  assign _T_3280 = {_T_3109,_T_3108,_T_3107,_T_3114,_T_3113,_T_3112,_T_3111,_T_3110}; // @[Mux.scala 19:72:@1605.4]
  assign _T_3282 = _T_2350 ? _T_3280 : 8'h0; // @[Mux.scala 19:72:@1606.4]
  assign _T_3289 = {_T_3148,_T_3147,_T_3154,_T_3153,_T_3152,_T_3151,_T_3150,_T_3149}; // @[Mux.scala 19:72:@1613.4]
  assign _T_3291 = _T_2351 ? _T_3289 : 8'h0; // @[Mux.scala 19:72:@1614.4]
  assign _T_3298 = {_T_3187,_T_3194,_T_3193,_T_3192,_T_3191,_T_3190,_T_3189,_T_3188}; // @[Mux.scala 19:72:@1621.4]
  assign _T_3300 = _T_2352 ? _T_3298 : 8'h0; // @[Mux.scala 19:72:@1622.4]
  assign _T_3301 = _T_3237 | _T_3246; // @[Mux.scala 19:72:@1623.4]
  assign _T_3302 = _T_3301 | _T_3255; // @[Mux.scala 19:72:@1624.4]
  assign _T_3303 = _T_3302 | _T_3264; // @[Mux.scala 19:72:@1625.4]
  assign _T_3304 = _T_3303 | _T_3273; // @[Mux.scala 19:72:@1626.4]
  assign _T_3305 = _T_3304 | _T_3282; // @[Mux.scala 19:72:@1627.4]
  assign _T_3306 = _T_3305 | _T_3291; // @[Mux.scala 19:72:@1628.4]
  assign _T_3307 = _T_3306 | _T_3300; // @[Mux.scala 19:72:@1629.4]
  assign inputDataPriorityPorts_0_0 = _T_3307[0]; // @[Mux.scala 19:72:@1633.4]
  assign inputDataPriorityPorts_0_1 = _T_3307[1]; // @[Mux.scala 19:72:@1635.4]
  assign inputDataPriorityPorts_0_2 = _T_3307[2]; // @[Mux.scala 19:72:@1637.4]
  assign inputDataPriorityPorts_0_3 = _T_3307[3]; // @[Mux.scala 19:72:@1639.4]
  assign inputDataPriorityPorts_0_4 = _T_3307[4]; // @[Mux.scala 19:72:@1641.4]
  assign inputDataPriorityPorts_0_5 = _T_3307[5]; // @[Mux.scala 19:72:@1643.4]
  assign inputDataPriorityPorts_0_6 = _T_3307[6]; // @[Mux.scala 19:72:@1645.4]
  assign inputDataPriorityPorts_0_7 = _T_3307[7]; // @[Mux.scala 19:72:@1647.4]
  assign _T_3389 = inputAddrPriorityPorts_0_0 & _T_2266; // @[StoreQueue.scala 209:52:@1663.6]
  assign _T_3390 = _T_3389 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@1664.6]
  assign _GEN_304 = _T_3390 ? io_addressFromStorePorts_0 : addrQ_0; // @[StoreQueue.scala 210:40:@1668.6]
  assign _GEN_305 = _T_3390 ? 1'h1 : addrKnown_0; // @[StoreQueue.scala 210:40:@1668.6]
  assign _T_3406 = inputDataPriorityPorts_0_0 & _T_2304; // @[StoreQueue.scala 215:52:@1673.6]
  assign _T_3407 = _T_3406 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@1674.6]
  assign _GEN_306 = _T_3407 ? io_dataFromStorePorts_0 : dataQ_0; // @[StoreQueue.scala 216:40:@1678.6]
  assign _GEN_307 = _T_3407 ? 1'h1 : dataKnown_0; // @[StoreQueue.scala 216:40:@1678.6]
  assign _GEN_308 = initBits_0 ? 1'h0 : _GEN_305; // @[StoreQueue.scala 204:35:@1657.4]
  assign _GEN_309 = initBits_0 ? 1'h0 : _GEN_307; // @[StoreQueue.scala 204:35:@1657.4]
  assign _GEN_310 = initBits_0 ? addrQ_0 : _GEN_304; // @[StoreQueue.scala 204:35:@1657.4]
  assign _GEN_311 = initBits_0 ? dataQ_0 : _GEN_306; // @[StoreQueue.scala 204:35:@1657.4]
  assign _T_3425 = inputAddrPriorityPorts_0_1 & _T_2269; // @[StoreQueue.scala 209:52:@1689.6]
  assign _T_3426 = _T_3425 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@1690.6]
  assign _GEN_312 = _T_3426 ? io_addressFromStorePorts_0 : addrQ_1; // @[StoreQueue.scala 210:40:@1694.6]
  assign _GEN_313 = _T_3426 ? 1'h1 : addrKnown_1; // @[StoreQueue.scala 210:40:@1694.6]
  assign _T_3442 = inputDataPriorityPorts_0_1 & _T_2307; // @[StoreQueue.scala 215:52:@1699.6]
  assign _T_3443 = _T_3442 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@1700.6]
  assign _GEN_314 = _T_3443 ? io_dataFromStorePorts_0 : dataQ_1; // @[StoreQueue.scala 216:40:@1704.6]
  assign _GEN_315 = _T_3443 ? 1'h1 : dataKnown_1; // @[StoreQueue.scala 216:40:@1704.6]
  assign _GEN_316 = initBits_1 ? 1'h0 : _GEN_313; // @[StoreQueue.scala 204:35:@1683.4]
  assign _GEN_317 = initBits_1 ? 1'h0 : _GEN_315; // @[StoreQueue.scala 204:35:@1683.4]
  assign _GEN_318 = initBits_1 ? addrQ_1 : _GEN_312; // @[StoreQueue.scala 204:35:@1683.4]
  assign _GEN_319 = initBits_1 ? dataQ_1 : _GEN_314; // @[StoreQueue.scala 204:35:@1683.4]
  assign _T_3461 = inputAddrPriorityPorts_0_2 & _T_2272; // @[StoreQueue.scala 209:52:@1715.6]
  assign _T_3462 = _T_3461 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@1716.6]
  assign _GEN_320 = _T_3462 ? io_addressFromStorePorts_0 : addrQ_2; // @[StoreQueue.scala 210:40:@1720.6]
  assign _GEN_321 = _T_3462 ? 1'h1 : addrKnown_2; // @[StoreQueue.scala 210:40:@1720.6]
  assign _T_3478 = inputDataPriorityPorts_0_2 & _T_2310; // @[StoreQueue.scala 215:52:@1725.6]
  assign _T_3479 = _T_3478 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@1726.6]
  assign _GEN_322 = _T_3479 ? io_dataFromStorePorts_0 : dataQ_2; // @[StoreQueue.scala 216:40:@1730.6]
  assign _GEN_323 = _T_3479 ? 1'h1 : dataKnown_2; // @[StoreQueue.scala 216:40:@1730.6]
  assign _GEN_324 = initBits_2 ? 1'h0 : _GEN_321; // @[StoreQueue.scala 204:35:@1709.4]
  assign _GEN_325 = initBits_2 ? 1'h0 : _GEN_323; // @[StoreQueue.scala 204:35:@1709.4]
  assign _GEN_326 = initBits_2 ? addrQ_2 : _GEN_320; // @[StoreQueue.scala 204:35:@1709.4]
  assign _GEN_327 = initBits_2 ? dataQ_2 : _GEN_322; // @[StoreQueue.scala 204:35:@1709.4]
  assign _T_3497 = inputAddrPriorityPorts_0_3 & _T_2275; // @[StoreQueue.scala 209:52:@1741.6]
  assign _T_3498 = _T_3497 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@1742.6]
  assign _GEN_328 = _T_3498 ? io_addressFromStorePorts_0 : addrQ_3; // @[StoreQueue.scala 210:40:@1746.6]
  assign _GEN_329 = _T_3498 ? 1'h1 : addrKnown_3; // @[StoreQueue.scala 210:40:@1746.6]
  assign _T_3514 = inputDataPriorityPorts_0_3 & _T_2313; // @[StoreQueue.scala 215:52:@1751.6]
  assign _T_3515 = _T_3514 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@1752.6]
  assign _GEN_330 = _T_3515 ? io_dataFromStorePorts_0 : dataQ_3; // @[StoreQueue.scala 216:40:@1756.6]
  assign _GEN_331 = _T_3515 ? 1'h1 : dataKnown_3; // @[StoreQueue.scala 216:40:@1756.6]
  assign _GEN_332 = initBits_3 ? 1'h0 : _GEN_329; // @[StoreQueue.scala 204:35:@1735.4]
  assign _GEN_333 = initBits_3 ? 1'h0 : _GEN_331; // @[StoreQueue.scala 204:35:@1735.4]
  assign _GEN_334 = initBits_3 ? addrQ_3 : _GEN_328; // @[StoreQueue.scala 204:35:@1735.4]
  assign _GEN_335 = initBits_3 ? dataQ_3 : _GEN_330; // @[StoreQueue.scala 204:35:@1735.4]
  assign _T_3533 = inputAddrPriorityPorts_0_4 & _T_2278; // @[StoreQueue.scala 209:52:@1767.6]
  assign _T_3534 = _T_3533 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@1768.6]
  assign _GEN_336 = _T_3534 ? io_addressFromStorePorts_0 : addrQ_4; // @[StoreQueue.scala 210:40:@1772.6]
  assign _GEN_337 = _T_3534 ? 1'h1 : addrKnown_4; // @[StoreQueue.scala 210:40:@1772.6]
  assign _T_3550 = inputDataPriorityPorts_0_4 & _T_2316; // @[StoreQueue.scala 215:52:@1777.6]
  assign _T_3551 = _T_3550 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@1778.6]
  assign _GEN_338 = _T_3551 ? io_dataFromStorePorts_0 : dataQ_4; // @[StoreQueue.scala 216:40:@1782.6]
  assign _GEN_339 = _T_3551 ? 1'h1 : dataKnown_4; // @[StoreQueue.scala 216:40:@1782.6]
  assign _GEN_340 = initBits_4 ? 1'h0 : _GEN_337; // @[StoreQueue.scala 204:35:@1761.4]
  assign _GEN_341 = initBits_4 ? 1'h0 : _GEN_339; // @[StoreQueue.scala 204:35:@1761.4]
  assign _GEN_342 = initBits_4 ? addrQ_4 : _GEN_336; // @[StoreQueue.scala 204:35:@1761.4]
  assign _GEN_343 = initBits_4 ? dataQ_4 : _GEN_338; // @[StoreQueue.scala 204:35:@1761.4]
  assign _T_3569 = inputAddrPriorityPorts_0_5 & _T_2281; // @[StoreQueue.scala 209:52:@1793.6]
  assign _T_3570 = _T_3569 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@1794.6]
  assign _GEN_344 = _T_3570 ? io_addressFromStorePorts_0 : addrQ_5; // @[StoreQueue.scala 210:40:@1798.6]
  assign _GEN_345 = _T_3570 ? 1'h1 : addrKnown_5; // @[StoreQueue.scala 210:40:@1798.6]
  assign _T_3586 = inputDataPriorityPorts_0_5 & _T_2319; // @[StoreQueue.scala 215:52:@1803.6]
  assign _T_3587 = _T_3586 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@1804.6]
  assign _GEN_346 = _T_3587 ? io_dataFromStorePorts_0 : dataQ_5; // @[StoreQueue.scala 216:40:@1808.6]
  assign _GEN_347 = _T_3587 ? 1'h1 : dataKnown_5; // @[StoreQueue.scala 216:40:@1808.6]
  assign _GEN_348 = initBits_5 ? 1'h0 : _GEN_345; // @[StoreQueue.scala 204:35:@1787.4]
  assign _GEN_349 = initBits_5 ? 1'h0 : _GEN_347; // @[StoreQueue.scala 204:35:@1787.4]
  assign _GEN_350 = initBits_5 ? addrQ_5 : _GEN_344; // @[StoreQueue.scala 204:35:@1787.4]
  assign _GEN_351 = initBits_5 ? dataQ_5 : _GEN_346; // @[StoreQueue.scala 204:35:@1787.4]
  assign _T_3605 = inputAddrPriorityPorts_0_6 & _T_2284; // @[StoreQueue.scala 209:52:@1819.6]
  assign _T_3606 = _T_3605 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@1820.6]
  assign _GEN_352 = _T_3606 ? io_addressFromStorePorts_0 : addrQ_6; // @[StoreQueue.scala 210:40:@1824.6]
  assign _GEN_353 = _T_3606 ? 1'h1 : addrKnown_6; // @[StoreQueue.scala 210:40:@1824.6]
  assign _T_3622 = inputDataPriorityPorts_0_6 & _T_2322; // @[StoreQueue.scala 215:52:@1829.6]
  assign _T_3623 = _T_3622 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@1830.6]
  assign _GEN_354 = _T_3623 ? io_dataFromStorePorts_0 : dataQ_6; // @[StoreQueue.scala 216:40:@1834.6]
  assign _GEN_355 = _T_3623 ? 1'h1 : dataKnown_6; // @[StoreQueue.scala 216:40:@1834.6]
  assign _GEN_356 = initBits_6 ? 1'h0 : _GEN_353; // @[StoreQueue.scala 204:35:@1813.4]
  assign _GEN_357 = initBits_6 ? 1'h0 : _GEN_355; // @[StoreQueue.scala 204:35:@1813.4]
  assign _GEN_358 = initBits_6 ? addrQ_6 : _GEN_352; // @[StoreQueue.scala 204:35:@1813.4]
  assign _GEN_359 = initBits_6 ? dataQ_6 : _GEN_354; // @[StoreQueue.scala 204:35:@1813.4]
  assign _T_3641 = inputAddrPriorityPorts_0_7 & _T_2287; // @[StoreQueue.scala 209:52:@1845.6]
  assign _T_3642 = _T_3641 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@1846.6]
  assign _GEN_360 = _T_3642 ? io_addressFromStorePorts_0 : addrQ_7; // @[StoreQueue.scala 210:40:@1850.6]
  assign _GEN_361 = _T_3642 ? 1'h1 : addrKnown_7; // @[StoreQueue.scala 210:40:@1850.6]
  assign _T_3658 = inputDataPriorityPorts_0_7 & _T_2325; // @[StoreQueue.scala 215:52:@1855.6]
  assign _T_3659 = _T_3658 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@1856.6]
  assign _GEN_362 = _T_3659 ? io_dataFromStorePorts_0 : dataQ_7; // @[StoreQueue.scala 216:40:@1860.6]
  assign _GEN_363 = _T_3659 ? 1'h1 : dataKnown_7; // @[StoreQueue.scala 216:40:@1860.6]
  assign _GEN_364 = initBits_7 ? 1'h0 : _GEN_361; // @[StoreQueue.scala 204:35:@1839.4]
  assign _GEN_365 = initBits_7 ? 1'h0 : _GEN_363; // @[StoreQueue.scala 204:35:@1839.4]
  assign _GEN_366 = initBits_7 ? addrQ_7 : _GEN_360; // @[StoreQueue.scala 204:35:@1839.4]
  assign _GEN_367 = initBits_7 ? dataQ_7 : _GEN_362; // @[StoreQueue.scala 204:35:@1839.4]
  assign _T_3673 = storeRequest & io_memIsReadyForStores; // @[StoreQueue.scala 229:23:@1865.4]
  assign _T_3676 = head + 3'h1; // @[util.scala 10:8:@1867.6]
  assign _GEN_32 = _T_3676 % 4'h8; // @[util.scala 10:14:@1868.6]
  assign _T_3677 = _GEN_32[3:0]; // @[util.scala 10:14:@1868.6]
  assign _GEN_368 = _T_3673 ? _T_3677 : {{1'd0}, head}; // @[StoreQueue.scala 229:50:@1866.4]
  assign _T_3679 = tail + io_bbNumStores; // @[util.scala 10:8:@1872.6]
  assign _GEN_33 = _T_3679 % 4'h8; // @[util.scala 10:14:@1873.6]
  assign _T_3680 = _GEN_33[3:0]; // @[util.scala 10:14:@1873.6]
  assign _GEN_369 = io_bbStart ? _T_3680 : {{1'd0}, tail}; // @[StoreQueue.scala 233:20:@1871.4]
  assign _T_3682 = allocatedEntries_0 == 1'h0; // @[StoreQueue.scala 237:84:@1876.4]
  assign _T_3683 = storeCompleted_0 | _T_3682; // @[StoreQueue.scala 237:81:@1877.4]
  assign _T_3685 = allocatedEntries_1 == 1'h0; // @[StoreQueue.scala 237:84:@1878.4]
  assign _T_3686 = storeCompleted_1 | _T_3685; // @[StoreQueue.scala 237:81:@1879.4]
  assign _T_3688 = allocatedEntries_2 == 1'h0; // @[StoreQueue.scala 237:84:@1880.4]
  assign _T_3689 = storeCompleted_2 | _T_3688; // @[StoreQueue.scala 237:81:@1881.4]
  assign _T_3691 = allocatedEntries_3 == 1'h0; // @[StoreQueue.scala 237:84:@1882.4]
  assign _T_3692 = storeCompleted_3 | _T_3691; // @[StoreQueue.scala 237:81:@1883.4]
  assign _T_3694 = allocatedEntries_4 == 1'h0; // @[StoreQueue.scala 237:84:@1884.4]
  assign _T_3695 = storeCompleted_4 | _T_3694; // @[StoreQueue.scala 237:81:@1885.4]
  assign _T_3697 = allocatedEntries_5 == 1'h0; // @[StoreQueue.scala 237:84:@1886.4]
  assign _T_3698 = storeCompleted_5 | _T_3697; // @[StoreQueue.scala 237:81:@1887.4]
  assign _T_3700 = allocatedEntries_6 == 1'h0; // @[StoreQueue.scala 237:84:@1888.4]
  assign _T_3701 = storeCompleted_6 | _T_3700; // @[StoreQueue.scala 237:81:@1889.4]
  assign _T_3703 = allocatedEntries_7 == 1'h0; // @[StoreQueue.scala 237:84:@1890.4]
  assign _T_3704 = storeCompleted_7 | _T_3703; // @[StoreQueue.scala 237:81:@1891.4]
  assign _T_3721 = _T_3683 & _T_3686; // @[StoreQueue.scala 237:98:@1902.4]
  assign _T_3722 = _T_3721 & _T_3689; // @[StoreQueue.scala 237:98:@1903.4]
  assign _T_3723 = _T_3722 & _T_3692; // @[StoreQueue.scala 237:98:@1904.4]
  assign _T_3724 = _T_3723 & _T_3695; // @[StoreQueue.scala 237:98:@1905.4]
  assign _T_3725 = _T_3724 & _T_3698; // @[StoreQueue.scala 237:98:@1906.4]
  assign _T_3726 = _T_3725 & _T_3701; // @[StoreQueue.scala 237:98:@1907.4]
  assign _GEN_371 = 3'h1 == head ? dataQ_1 : dataQ_0; // @[StoreQueue.scala 252:21:@1945.4]
  assign _GEN_372 = 3'h2 == head ? dataQ_2 : _GEN_371; // @[StoreQueue.scala 252:21:@1945.4]
  assign _GEN_373 = 3'h3 == head ? dataQ_3 : _GEN_372; // @[StoreQueue.scala 252:21:@1945.4]
  assign _GEN_374 = 3'h4 == head ? dataQ_4 : _GEN_373; // @[StoreQueue.scala 252:21:@1945.4]
  assign _GEN_375 = 3'h5 == head ? dataQ_5 : _GEN_374; // @[StoreQueue.scala 252:21:@1945.4]
  assign _GEN_376 = 3'h6 == head ? dataQ_6 : _GEN_375; // @[StoreQueue.scala 252:21:@1945.4]
  assign io_storeTail = tail; // @[StoreQueue.scala 246:16:@1911.4]
  assign io_storeHead = head; // @[StoreQueue.scala 245:16:@1910.4]
  assign io_storeEmpty = _T_3726 & _T_3704; // @[StoreQueue.scala 237:17:@1909.4]
  assign io_storeAddrDone_0 = addrKnown_0; // @[StoreQueue.scala 250:20:@1936.4]
  assign io_storeAddrDone_1 = addrKnown_1; // @[StoreQueue.scala 250:20:@1937.4]
  assign io_storeAddrDone_2 = addrKnown_2; // @[StoreQueue.scala 250:20:@1938.4]
  assign io_storeAddrDone_3 = addrKnown_3; // @[StoreQueue.scala 250:20:@1939.4]
  assign io_storeAddrDone_4 = addrKnown_4; // @[StoreQueue.scala 250:20:@1940.4]
  assign io_storeAddrDone_5 = addrKnown_5; // @[StoreQueue.scala 250:20:@1941.4]
  assign io_storeAddrDone_6 = addrKnown_6; // @[StoreQueue.scala 250:20:@1942.4]
  assign io_storeAddrDone_7 = addrKnown_7; // @[StoreQueue.scala 250:20:@1943.4]
  assign io_storeDataDone_0 = dataKnown_0; // @[StoreQueue.scala 249:20:@1928.4]
  assign io_storeDataDone_1 = dataKnown_1; // @[StoreQueue.scala 249:20:@1929.4]
  assign io_storeDataDone_2 = dataKnown_2; // @[StoreQueue.scala 249:20:@1930.4]
  assign io_storeDataDone_3 = dataKnown_3; // @[StoreQueue.scala 249:20:@1931.4]
  assign io_storeDataDone_4 = dataKnown_4; // @[StoreQueue.scala 249:20:@1932.4]
  assign io_storeDataDone_5 = dataKnown_5; // @[StoreQueue.scala 249:20:@1933.4]
  assign io_storeDataDone_6 = dataKnown_6; // @[StoreQueue.scala 249:20:@1934.4]
  assign io_storeDataDone_7 = dataKnown_7; // @[StoreQueue.scala 249:20:@1935.4]
  assign io_storeAddrQueue_0 = addrQ_0; // @[StoreQueue.scala 247:21:@1912.4]
  assign io_storeAddrQueue_1 = addrQ_1; // @[StoreQueue.scala 247:21:@1913.4]
  assign io_storeAddrQueue_2 = addrQ_2; // @[StoreQueue.scala 247:21:@1914.4]
  assign io_storeAddrQueue_3 = addrQ_3; // @[StoreQueue.scala 247:21:@1915.4]
  assign io_storeAddrQueue_4 = addrQ_4; // @[StoreQueue.scala 247:21:@1916.4]
  assign io_storeAddrQueue_5 = addrQ_5; // @[StoreQueue.scala 247:21:@1917.4]
  assign io_storeAddrQueue_6 = addrQ_6; // @[StoreQueue.scala 247:21:@1918.4]
  assign io_storeAddrQueue_7 = addrQ_7; // @[StoreQueue.scala 247:21:@1919.4]
  assign io_storeDataQueue_0 = dataQ_0; // @[StoreQueue.scala 248:21:@1920.4]
  assign io_storeDataQueue_1 = dataQ_1; // @[StoreQueue.scala 248:21:@1921.4]
  assign io_storeDataQueue_2 = dataQ_2; // @[StoreQueue.scala 248:21:@1922.4]
  assign io_storeDataQueue_3 = dataQ_3; // @[StoreQueue.scala 248:21:@1923.4]
  assign io_storeDataQueue_4 = dataQ_4; // @[StoreQueue.scala 248:21:@1924.4]
  assign io_storeDataQueue_5 = dataQ_5; // @[StoreQueue.scala 248:21:@1925.4]
  assign io_storeDataQueue_6 = dataQ_6; // @[StoreQueue.scala 248:21:@1926.4]
  assign io_storeDataQueue_7 = dataQ_7; // @[StoreQueue.scala 248:21:@1927.4]
  assign io_storeAddrToMem = 3'h7 == head ? addrQ_7 : _GEN_262; // @[StoreQueue.scala 253:21:@1946.4]
  assign io_storeDataToMem = 3'h7 == head ? dataQ_7 : _GEN_376; // @[StoreQueue.scala 252:21:@1945.4]
  assign io_storeEnableToMem = _T_1933 & _T_1942; // @[StoreQueue.scala 251:23:@1944.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  portQ_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  portQ_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  portQ_2 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  portQ_3 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  portQ_4 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  portQ_5 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  portQ_6 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  portQ_7 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  addrQ_0 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  addrQ_1 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  addrQ_2 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  addrQ_3 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  addrQ_4 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  addrQ_5 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  addrQ_6 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  addrQ_7 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  dataQ_0 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  dataQ_1 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  dataQ_2 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  dataQ_3 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  dataQ_4 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  dataQ_5 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  dataQ_6 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  dataQ_7 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrKnown_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrKnown_1 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrKnown_2 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrKnown_3 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrKnown_4 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrKnown_5 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrKnown_6 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrKnown_7 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  dataKnown_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  dataKnown_1 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  dataKnown_2 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  dataKnown_3 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  dataKnown_4 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  dataKnown_5 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  dataKnown_6 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  dataKnown_7 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  storeCompleted_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  storeCompleted_1 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  storeCompleted_2 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  storeCompleted_3 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  storeCompleted_4 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  storeCompleted_5 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  storeCompleted_6 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  storeCompleted_7 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  checkBits_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  checkBits_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  checkBits_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  checkBits_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  checkBits_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  checkBits_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  checkBits_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  checkBits_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  previousLoadHead = _RAND_74[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 3'h0;
    end else begin
      head <= _GEN_368[2:0];
    end
    if (reset) begin
      tail <= 3'h0;
    end else begin
      tail <= _GEN_369[2:0];
    end
    if (reset) begin
      offsetQ_0 <= 3'h0;
    end else begin
      if (initBits_0) begin
        if (3'h7 == _T_1060) begin
          offsetQ_0 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1060) begin
            offsetQ_0 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1060) begin
              offsetQ_0 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1060) begin
                offsetQ_0 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1060) begin
                  offsetQ_0 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1060) begin
                    offsetQ_0 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1060) begin
                      offsetQ_0 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_0 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 3'h0;
    end else begin
      if (initBits_1) begin
        if (3'h7 == _T_1078) begin
          offsetQ_1 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1078) begin
            offsetQ_1 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1078) begin
              offsetQ_1 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1078) begin
                offsetQ_1 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1078) begin
                  offsetQ_1 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1078) begin
                    offsetQ_1 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1078) begin
                      offsetQ_1 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_1 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 3'h0;
    end else begin
      if (initBits_2) begin
        if (3'h7 == _T_1096) begin
          offsetQ_2 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1096) begin
            offsetQ_2 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1096) begin
              offsetQ_2 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1096) begin
                offsetQ_2 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1096) begin
                  offsetQ_2 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1096) begin
                    offsetQ_2 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1096) begin
                      offsetQ_2 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_2 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 3'h0;
    end else begin
      if (initBits_3) begin
        if (3'h7 == _T_1114) begin
          offsetQ_3 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1114) begin
            offsetQ_3 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1114) begin
              offsetQ_3 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1114) begin
                offsetQ_3 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1114) begin
                  offsetQ_3 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1114) begin
                    offsetQ_3 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1114) begin
                      offsetQ_3 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_3 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 3'h0;
    end else begin
      if (initBits_4) begin
        if (3'h7 == _T_1132) begin
          offsetQ_4 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1132) begin
            offsetQ_4 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1132) begin
              offsetQ_4 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1132) begin
                offsetQ_4 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1132) begin
                  offsetQ_4 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1132) begin
                    offsetQ_4 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1132) begin
                      offsetQ_4 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_4 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 3'h0;
    end else begin
      if (initBits_5) begin
        if (3'h7 == _T_1150) begin
          offsetQ_5 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1150) begin
            offsetQ_5 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1150) begin
              offsetQ_5 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1150) begin
                offsetQ_5 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1150) begin
                  offsetQ_5 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1150) begin
                    offsetQ_5 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1150) begin
                      offsetQ_5 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_5 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 3'h0;
    end else begin
      if (initBits_6) begin
        if (3'h7 == _T_1168) begin
          offsetQ_6 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1168) begin
            offsetQ_6 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1168) begin
              offsetQ_6 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1168) begin
                offsetQ_6 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1168) begin
                  offsetQ_6 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1168) begin
                    offsetQ_6 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1168) begin
                      offsetQ_6 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_6 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 3'h0;
    end else begin
      if (initBits_7) begin
        if (3'h7 == _T_1186) begin
          offsetQ_7 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1186) begin
            offsetQ_7 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1186) begin
              offsetQ_7 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1186) begin
                offsetQ_7 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1186) begin
                  offsetQ_7 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1186) begin
                    offsetQ_7 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1186) begin
                      offsetQ_7 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_7 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        portQ_0 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        portQ_1 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        portQ_2 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        portQ_3 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        portQ_4 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        portQ_5 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        portQ_6 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        portQ_7 <= 1'h0;
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_3390) begin
          addrQ_0 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_3426) begin
          addrQ_1 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_3462) begin
          addrQ_2 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_3498) begin
          addrQ_3 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_3534) begin
          addrQ_4 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_3570) begin
          addrQ_5 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_3606) begin
          addrQ_6 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_3642) begin
          addrQ_7 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_3407) begin
          dataQ_0 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_3443) begin
          dataQ_1 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_3479) begin
          dataQ_2 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_3515) begin
          dataQ_3 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_3551) begin
          dataQ_4 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_3587) begin
          dataQ_5 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_3623) begin
          dataQ_6 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_3659) begin
          dataQ_7 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_3390) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_3426) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_3462) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_3498) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_3534) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_3570) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_3606) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_3642) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_3407) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_3443) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_3479) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_3515) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_3551) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_3587) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_3623) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_3659) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1030;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1031;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1032;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1033;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1034;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1035;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1036;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1037;
    end
    if (reset) begin
      storeCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        storeCompleted_0 <= 1'h0;
      end else begin
        if (_T_1947) begin
          storeCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        storeCompleted_1 <= 1'h0;
      end else begin
        if (_T_1953) begin
          storeCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        storeCompleted_2 <= 1'h0;
      end else begin
        if (_T_1959) begin
          storeCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        storeCompleted_3 <= 1'h0;
      end else begin
        if (_T_1965) begin
          storeCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        storeCompleted_4 <= 1'h0;
      end else begin
        if (_T_1971) begin
          storeCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        storeCompleted_5 <= 1'h0;
      end else begin
        if (_T_1977) begin
          storeCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        storeCompleted_6 <= 1'h0;
      end else begin
        if (_T_1983) begin
          storeCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        storeCompleted_7 <= 1'h0;
      end else begin
        if (_T_1989) begin
          storeCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_1213;
      end else begin
        if (io_loadEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_1217) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_1225) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_1243;
      end else begin
        if (io_loadEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_1247) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_1255) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_1273;
      end else begin
        if (io_loadEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_1277) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_1285) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_1303;
      end else begin
        if (io_loadEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_1307) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_1315) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_1333;
      end else begin
        if (io_loadEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_1337) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_1345) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_1363;
      end else begin
        if (io_loadEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_1367) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_1375) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_1393;
      end else begin
        if (io_loadEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_1397) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_1405) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_1423;
      end else begin
        if (io_loadEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_1427) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_1435) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    previousLoadHead <= io_loadHead;
  end
endmodule
module LOAD_QUEUE_LSQ_dist( // @[:@1948.2]
  input         clock, // @[:@1949.4]
  input         reset, // @[:@1950.4]
  input         io_bbStart, // @[:@1951.4]
  input  [2:0]  io_bbLoadOffsets_0, // @[:@1951.4]
  input  [2:0]  io_bbLoadOffsets_1, // @[:@1951.4]
  input  [2:0]  io_bbLoadOffsets_2, // @[:@1951.4]
  input  [2:0]  io_bbLoadOffsets_3, // @[:@1951.4]
  input  [2:0]  io_bbLoadOffsets_4, // @[:@1951.4]
  input  [2:0]  io_bbLoadOffsets_5, // @[:@1951.4]
  input  [2:0]  io_bbLoadOffsets_6, // @[:@1951.4]
  input  [2:0]  io_bbLoadOffsets_7, // @[:@1951.4]
  input  [2:0]  io_bbLoadPorts_0, // @[:@1951.4]
  input  [2:0]  io_bbLoadPorts_1, // @[:@1951.4]
  input  [2:0]  io_bbLoadPorts_2, // @[:@1951.4]
  input  [2:0]  io_bbNumLoads, // @[:@1951.4]
  output [2:0]  io_loadTail, // @[:@1951.4]
  output [2:0]  io_loadHead, // @[:@1951.4]
  output        io_loadEmpty, // @[:@1951.4]
  input  [2:0]  io_storeTail, // @[:@1951.4]
  input  [2:0]  io_storeHead, // @[:@1951.4]
  input         io_storeEmpty, // @[:@1951.4]
  input         io_storeAddrDone_0, // @[:@1951.4]
  input         io_storeAddrDone_1, // @[:@1951.4]
  input         io_storeAddrDone_2, // @[:@1951.4]
  input         io_storeAddrDone_3, // @[:@1951.4]
  input         io_storeAddrDone_4, // @[:@1951.4]
  input         io_storeAddrDone_5, // @[:@1951.4]
  input         io_storeAddrDone_6, // @[:@1951.4]
  input         io_storeAddrDone_7, // @[:@1951.4]
  input         io_storeDataDone_0, // @[:@1951.4]
  input         io_storeDataDone_1, // @[:@1951.4]
  input         io_storeDataDone_2, // @[:@1951.4]
  input         io_storeDataDone_3, // @[:@1951.4]
  input         io_storeDataDone_4, // @[:@1951.4]
  input         io_storeDataDone_5, // @[:@1951.4]
  input         io_storeDataDone_6, // @[:@1951.4]
  input         io_storeDataDone_7, // @[:@1951.4]
  input  [31:0] io_storeAddrQueue_0, // @[:@1951.4]
  input  [31:0] io_storeAddrQueue_1, // @[:@1951.4]
  input  [31:0] io_storeAddrQueue_2, // @[:@1951.4]
  input  [31:0] io_storeAddrQueue_3, // @[:@1951.4]
  input  [31:0] io_storeAddrQueue_4, // @[:@1951.4]
  input  [31:0] io_storeAddrQueue_5, // @[:@1951.4]
  input  [31:0] io_storeAddrQueue_6, // @[:@1951.4]
  input  [31:0] io_storeAddrQueue_7, // @[:@1951.4]
  input  [31:0] io_storeDataQueue_0, // @[:@1951.4]
  input  [31:0] io_storeDataQueue_1, // @[:@1951.4]
  input  [31:0] io_storeDataQueue_2, // @[:@1951.4]
  input  [31:0] io_storeDataQueue_3, // @[:@1951.4]
  input  [31:0] io_storeDataQueue_4, // @[:@1951.4]
  input  [31:0] io_storeDataQueue_5, // @[:@1951.4]
  input  [31:0] io_storeDataQueue_6, // @[:@1951.4]
  input  [31:0] io_storeDataQueue_7, // @[:@1951.4]
  output        io_loadAddrDone_0, // @[:@1951.4]
  output        io_loadAddrDone_1, // @[:@1951.4]
  output        io_loadAddrDone_2, // @[:@1951.4]
  output        io_loadAddrDone_3, // @[:@1951.4]
  output        io_loadAddrDone_4, // @[:@1951.4]
  output        io_loadAddrDone_5, // @[:@1951.4]
  output        io_loadAddrDone_6, // @[:@1951.4]
  output        io_loadAddrDone_7, // @[:@1951.4]
  output        io_loadDataDone_0, // @[:@1951.4]
  output        io_loadDataDone_1, // @[:@1951.4]
  output        io_loadDataDone_2, // @[:@1951.4]
  output        io_loadDataDone_3, // @[:@1951.4]
  output        io_loadDataDone_4, // @[:@1951.4]
  output        io_loadDataDone_5, // @[:@1951.4]
  output        io_loadDataDone_6, // @[:@1951.4]
  output        io_loadDataDone_7, // @[:@1951.4]
  output [31:0] io_loadAddrQueue_0, // @[:@1951.4]
  output [31:0] io_loadAddrQueue_1, // @[:@1951.4]
  output [31:0] io_loadAddrQueue_2, // @[:@1951.4]
  output [31:0] io_loadAddrQueue_3, // @[:@1951.4]
  output [31:0] io_loadAddrQueue_4, // @[:@1951.4]
  output [31:0] io_loadAddrQueue_5, // @[:@1951.4]
  output [31:0] io_loadAddrQueue_6, // @[:@1951.4]
  output [31:0] io_loadAddrQueue_7, // @[:@1951.4]
  input         io_loadAddrEnable_0, // @[:@1951.4]
  input         io_loadAddrEnable_1, // @[:@1951.4]
  input         io_loadAddrEnable_2, // @[:@1951.4]
  input         io_loadAddrEnable_3, // @[:@1951.4]
  input         io_loadAddrEnable_4, // @[:@1951.4]
  input  [31:0] io_addrFromLoadPorts_0, // @[:@1951.4]
  input  [31:0] io_addrFromLoadPorts_1, // @[:@1951.4]
  input  [31:0] io_addrFromLoadPorts_2, // @[:@1951.4]
  input  [31:0] io_addrFromLoadPorts_3, // @[:@1951.4]
  input  [31:0] io_addrFromLoadPorts_4, // @[:@1951.4]
  input         io_loadPorts_0_ready, // @[:@1951.4]
  output        io_loadPorts_0_valid, // @[:@1951.4]
  output [31:0] io_loadPorts_0_bits, // @[:@1951.4]
  input         io_loadPorts_1_ready, // @[:@1951.4]
  output        io_loadPorts_1_valid, // @[:@1951.4]
  output [31:0] io_loadPorts_1_bits, // @[:@1951.4]
  input         io_loadPorts_2_ready, // @[:@1951.4]
  output        io_loadPorts_2_valid, // @[:@1951.4]
  output [31:0] io_loadPorts_2_bits, // @[:@1951.4]
  input         io_loadPorts_3_ready, // @[:@1951.4]
  output        io_loadPorts_3_valid, // @[:@1951.4]
  output [31:0] io_loadPorts_3_bits, // @[:@1951.4]
  input         io_loadPorts_4_ready, // @[:@1951.4]
  output        io_loadPorts_4_valid, // @[:@1951.4]
  output [31:0] io_loadPorts_4_bits, // @[:@1951.4]
  input  [31:0] io_loadDataFromMem, // @[:@1951.4]
  output [31:0] io_loadAddrToMem, // @[:@1951.4]
  output        io_loadEnableToMem, // @[:@1951.4]
  input         io_memIsReadyForLoads // @[:@1951.4]
);
  reg [2:0] head; // @[LoadQueue.scala 50:21:@1953.4]
  reg [31:0] _RAND_0;
  reg [2:0] tail; // @[LoadQueue.scala 51:21:@1954.4]
  reg [31:0] _RAND_1;
  reg [2:0] offsetQ_0; // @[LoadQueue.scala 53:24:@1964.4]
  reg [31:0] _RAND_2;
  reg [2:0] offsetQ_1; // @[LoadQueue.scala 53:24:@1964.4]
  reg [31:0] _RAND_3;
  reg [2:0] offsetQ_2; // @[LoadQueue.scala 53:24:@1964.4]
  reg [31:0] _RAND_4;
  reg [2:0] offsetQ_3; // @[LoadQueue.scala 53:24:@1964.4]
  reg [31:0] _RAND_5;
  reg [2:0] offsetQ_4; // @[LoadQueue.scala 53:24:@1964.4]
  reg [31:0] _RAND_6;
  reg [2:0] offsetQ_5; // @[LoadQueue.scala 53:24:@1964.4]
  reg [31:0] _RAND_7;
  reg [2:0] offsetQ_6; // @[LoadQueue.scala 53:24:@1964.4]
  reg [31:0] _RAND_8;
  reg [2:0] offsetQ_7; // @[LoadQueue.scala 53:24:@1964.4]
  reg [31:0] _RAND_9;
  reg [2:0] portQ_0; // @[LoadQueue.scala 54:22:@1974.4]
  reg [31:0] _RAND_10;
  reg [2:0] portQ_1; // @[LoadQueue.scala 54:22:@1974.4]
  reg [31:0] _RAND_11;
  reg [2:0] portQ_2; // @[LoadQueue.scala 54:22:@1974.4]
  reg [31:0] _RAND_12;
  reg [2:0] portQ_3; // @[LoadQueue.scala 54:22:@1974.4]
  reg [31:0] _RAND_13;
  reg [2:0] portQ_4; // @[LoadQueue.scala 54:22:@1974.4]
  reg [31:0] _RAND_14;
  reg [2:0] portQ_5; // @[LoadQueue.scala 54:22:@1974.4]
  reg [31:0] _RAND_15;
  reg [2:0] portQ_6; // @[LoadQueue.scala 54:22:@1974.4]
  reg [31:0] _RAND_16;
  reg [2:0] portQ_7; // @[LoadQueue.scala 54:22:@1974.4]
  reg [31:0] _RAND_17;
  reg [31:0] addrQ_0; // @[LoadQueue.scala 55:22:@1984.4]
  reg [31:0] _RAND_18;
  reg [31:0] addrQ_1; // @[LoadQueue.scala 55:22:@1984.4]
  reg [31:0] _RAND_19;
  reg [31:0] addrQ_2; // @[LoadQueue.scala 55:22:@1984.4]
  reg [31:0] _RAND_20;
  reg [31:0] addrQ_3; // @[LoadQueue.scala 55:22:@1984.4]
  reg [31:0] _RAND_21;
  reg [31:0] addrQ_4; // @[LoadQueue.scala 55:22:@1984.4]
  reg [31:0] _RAND_22;
  reg [31:0] addrQ_5; // @[LoadQueue.scala 55:22:@1984.4]
  reg [31:0] _RAND_23;
  reg [31:0] addrQ_6; // @[LoadQueue.scala 55:22:@1984.4]
  reg [31:0] _RAND_24;
  reg [31:0] addrQ_7; // @[LoadQueue.scala 55:22:@1984.4]
  reg [31:0] _RAND_25;
  reg [31:0] dataQ_0; // @[LoadQueue.scala 56:22:@1994.4]
  reg [31:0] _RAND_26;
  reg [31:0] dataQ_1; // @[LoadQueue.scala 56:22:@1994.4]
  reg [31:0] _RAND_27;
  reg [31:0] dataQ_2; // @[LoadQueue.scala 56:22:@1994.4]
  reg [31:0] _RAND_28;
  reg [31:0] dataQ_3; // @[LoadQueue.scala 56:22:@1994.4]
  reg [31:0] _RAND_29;
  reg [31:0] dataQ_4; // @[LoadQueue.scala 56:22:@1994.4]
  reg [31:0] _RAND_30;
  reg [31:0] dataQ_5; // @[LoadQueue.scala 56:22:@1994.4]
  reg [31:0] _RAND_31;
  reg [31:0] dataQ_6; // @[LoadQueue.scala 56:22:@1994.4]
  reg [31:0] _RAND_32;
  reg [31:0] dataQ_7; // @[LoadQueue.scala 56:22:@1994.4]
  reg [31:0] _RAND_33;
  reg  addrKnown_0; // @[LoadQueue.scala 57:26:@2004.4]
  reg [31:0] _RAND_34;
  reg  addrKnown_1; // @[LoadQueue.scala 57:26:@2004.4]
  reg [31:0] _RAND_35;
  reg  addrKnown_2; // @[LoadQueue.scala 57:26:@2004.4]
  reg [31:0] _RAND_36;
  reg  addrKnown_3; // @[LoadQueue.scala 57:26:@2004.4]
  reg [31:0] _RAND_37;
  reg  addrKnown_4; // @[LoadQueue.scala 57:26:@2004.4]
  reg [31:0] _RAND_38;
  reg  addrKnown_5; // @[LoadQueue.scala 57:26:@2004.4]
  reg [31:0] _RAND_39;
  reg  addrKnown_6; // @[LoadQueue.scala 57:26:@2004.4]
  reg [31:0] _RAND_40;
  reg  addrKnown_7; // @[LoadQueue.scala 57:26:@2004.4]
  reg [31:0] _RAND_41;
  reg  dataKnown_0; // @[LoadQueue.scala 58:26:@2014.4]
  reg [31:0] _RAND_42;
  reg  dataKnown_1; // @[LoadQueue.scala 58:26:@2014.4]
  reg [31:0] _RAND_43;
  reg  dataKnown_2; // @[LoadQueue.scala 58:26:@2014.4]
  reg [31:0] _RAND_44;
  reg  dataKnown_3; // @[LoadQueue.scala 58:26:@2014.4]
  reg [31:0] _RAND_45;
  reg  dataKnown_4; // @[LoadQueue.scala 58:26:@2014.4]
  reg [31:0] _RAND_46;
  reg  dataKnown_5; // @[LoadQueue.scala 58:26:@2014.4]
  reg [31:0] _RAND_47;
  reg  dataKnown_6; // @[LoadQueue.scala 58:26:@2014.4]
  reg [31:0] _RAND_48;
  reg  dataKnown_7; // @[LoadQueue.scala 58:26:@2014.4]
  reg [31:0] _RAND_49;
  reg  loadCompleted_0; // @[LoadQueue.scala 59:30:@2024.4]
  reg [31:0] _RAND_50;
  reg  loadCompleted_1; // @[LoadQueue.scala 59:30:@2024.4]
  reg [31:0] _RAND_51;
  reg  loadCompleted_2; // @[LoadQueue.scala 59:30:@2024.4]
  reg [31:0] _RAND_52;
  reg  loadCompleted_3; // @[LoadQueue.scala 59:30:@2024.4]
  reg [31:0] _RAND_53;
  reg  loadCompleted_4; // @[LoadQueue.scala 59:30:@2024.4]
  reg [31:0] _RAND_54;
  reg  loadCompleted_5; // @[LoadQueue.scala 59:30:@2024.4]
  reg [31:0] _RAND_55;
  reg  loadCompleted_6; // @[LoadQueue.scala 59:30:@2024.4]
  reg [31:0] _RAND_56;
  reg  loadCompleted_7; // @[LoadQueue.scala 59:30:@2024.4]
  reg [31:0] _RAND_57;
  reg  allocatedEntries_0; // @[LoadQueue.scala 60:33:@2034.4]
  reg [31:0] _RAND_58;
  reg  allocatedEntries_1; // @[LoadQueue.scala 60:33:@2034.4]
  reg [31:0] _RAND_59;
  reg  allocatedEntries_2; // @[LoadQueue.scala 60:33:@2034.4]
  reg [31:0] _RAND_60;
  reg  allocatedEntries_3; // @[LoadQueue.scala 60:33:@2034.4]
  reg [31:0] _RAND_61;
  reg  allocatedEntries_4; // @[LoadQueue.scala 60:33:@2034.4]
  reg [31:0] _RAND_62;
  reg  allocatedEntries_5; // @[LoadQueue.scala 60:33:@2034.4]
  reg [31:0] _RAND_63;
  reg  allocatedEntries_6; // @[LoadQueue.scala 60:33:@2034.4]
  reg [31:0] _RAND_64;
  reg  allocatedEntries_7; // @[LoadQueue.scala 60:33:@2034.4]
  reg [31:0] _RAND_65;
  reg  bypassInitiated_0; // @[LoadQueue.scala 61:32:@2044.4]
  reg [31:0] _RAND_66;
  reg  bypassInitiated_1; // @[LoadQueue.scala 61:32:@2044.4]
  reg [31:0] _RAND_67;
  reg  bypassInitiated_2; // @[LoadQueue.scala 61:32:@2044.4]
  reg [31:0] _RAND_68;
  reg  bypassInitiated_3; // @[LoadQueue.scala 61:32:@2044.4]
  reg [31:0] _RAND_69;
  reg  bypassInitiated_4; // @[LoadQueue.scala 61:32:@2044.4]
  reg [31:0] _RAND_70;
  reg  bypassInitiated_5; // @[LoadQueue.scala 61:32:@2044.4]
  reg [31:0] _RAND_71;
  reg  bypassInitiated_6; // @[LoadQueue.scala 61:32:@2044.4]
  reg [31:0] _RAND_72;
  reg  bypassInitiated_7; // @[LoadQueue.scala 61:32:@2044.4]
  reg [31:0] _RAND_73;
  reg  checkBits_0; // @[LoadQueue.scala 62:26:@2054.4]
  reg [31:0] _RAND_74;
  reg  checkBits_1; // @[LoadQueue.scala 62:26:@2054.4]
  reg [31:0] _RAND_75;
  reg  checkBits_2; // @[LoadQueue.scala 62:26:@2054.4]
  reg [31:0] _RAND_76;
  reg  checkBits_3; // @[LoadQueue.scala 62:26:@2054.4]
  reg [31:0] _RAND_77;
  reg  checkBits_4; // @[LoadQueue.scala 62:26:@2054.4]
  reg [31:0] _RAND_78;
  reg  checkBits_5; // @[LoadQueue.scala 62:26:@2054.4]
  reg [31:0] _RAND_79;
  reg  checkBits_6; // @[LoadQueue.scala 62:26:@2054.4]
  reg [31:0] _RAND_80;
  reg  checkBits_7; // @[LoadQueue.scala 62:26:@2054.4]
  reg [31:0] _RAND_81;
  wire [4:0] _GEN_766; // @[util.scala 14:20:@2056.4]
  wire [5:0] _T_1044; // @[util.scala 14:20:@2056.4]
  wire [5:0] _T_1045; // @[util.scala 14:20:@2057.4]
  wire [4:0] _T_1046; // @[util.scala 14:20:@2058.4]
  wire [4:0] _GEN_0; // @[util.scala 14:25:@2059.4]
  wire [3:0] _T_1047; // @[util.scala 14:25:@2059.4]
  wire [3:0] _GEN_767; // @[LoadQueue.scala 71:46:@2060.4]
  wire  _T_1048; // @[LoadQueue.scala 71:46:@2060.4]
  wire  initBits_0; // @[LoadQueue.scala 71:63:@2061.4]
  wire [5:0] _T_1053; // @[util.scala 14:20:@2063.4]
  wire [5:0] _T_1054; // @[util.scala 14:20:@2064.4]
  wire [4:0] _T_1055; // @[util.scala 14:20:@2065.4]
  wire [4:0] _GEN_8; // @[util.scala 14:25:@2066.4]
  wire [3:0] _T_1056; // @[util.scala 14:25:@2066.4]
  wire  _T_1057; // @[LoadQueue.scala 71:46:@2067.4]
  wire  initBits_1; // @[LoadQueue.scala 71:63:@2068.4]
  wire [5:0] _T_1062; // @[util.scala 14:20:@2070.4]
  wire [5:0] _T_1063; // @[util.scala 14:20:@2071.4]
  wire [4:0] _T_1064; // @[util.scala 14:20:@2072.4]
  wire [4:0] _GEN_18; // @[util.scala 14:25:@2073.4]
  wire [3:0] _T_1065; // @[util.scala 14:25:@2073.4]
  wire  _T_1066; // @[LoadQueue.scala 71:46:@2074.4]
  wire  initBits_2; // @[LoadQueue.scala 71:63:@2075.4]
  wire [5:0] _T_1071; // @[util.scala 14:20:@2077.4]
  wire [5:0] _T_1072; // @[util.scala 14:20:@2078.4]
  wire [4:0] _T_1073; // @[util.scala 14:20:@2079.4]
  wire [4:0] _GEN_26; // @[util.scala 14:25:@2080.4]
  wire [3:0] _T_1074; // @[util.scala 14:25:@2080.4]
  wire  _T_1075; // @[LoadQueue.scala 71:46:@2081.4]
  wire  initBits_3; // @[LoadQueue.scala 71:63:@2082.4]
  wire [5:0] _T_1080; // @[util.scala 14:20:@2084.4]
  wire [5:0] _T_1081; // @[util.scala 14:20:@2085.4]
  wire [4:0] _T_1082; // @[util.scala 14:20:@2086.4]
  wire [4:0] _GEN_36; // @[util.scala 14:25:@2087.4]
  wire [3:0] _T_1083; // @[util.scala 14:25:@2087.4]
  wire  _T_1084; // @[LoadQueue.scala 71:46:@2088.4]
  wire  initBits_4; // @[LoadQueue.scala 71:63:@2089.4]
  wire [5:0] _T_1089; // @[util.scala 14:20:@2091.4]
  wire [5:0] _T_1090; // @[util.scala 14:20:@2092.4]
  wire [4:0] _T_1091; // @[util.scala 14:20:@2093.4]
  wire [4:0] _GEN_44; // @[util.scala 14:25:@2094.4]
  wire [3:0] _T_1092; // @[util.scala 14:25:@2094.4]
  wire  _T_1093; // @[LoadQueue.scala 71:46:@2095.4]
  wire  initBits_5; // @[LoadQueue.scala 71:63:@2096.4]
  wire [5:0] _T_1098; // @[util.scala 14:20:@2098.4]
  wire [5:0] _T_1099; // @[util.scala 14:20:@2099.4]
  wire [4:0] _T_1100; // @[util.scala 14:20:@2100.4]
  wire [4:0] _GEN_54; // @[util.scala 14:25:@2101.4]
  wire [3:0] _T_1101; // @[util.scala 14:25:@2101.4]
  wire  _T_1102; // @[LoadQueue.scala 71:46:@2102.4]
  wire  initBits_6; // @[LoadQueue.scala 71:63:@2103.4]
  wire [5:0] _T_1107; // @[util.scala 14:20:@2105.4]
  wire [5:0] _T_1108; // @[util.scala 14:20:@2106.4]
  wire [4:0] _T_1109; // @[util.scala 14:20:@2107.4]
  wire [4:0] _GEN_62; // @[util.scala 14:25:@2108.4]
  wire [3:0] _T_1110; // @[util.scala 14:25:@2108.4]
  wire  _T_1111; // @[LoadQueue.scala 71:46:@2109.4]
  wire  initBits_7; // @[LoadQueue.scala 71:63:@2110.4]
  wire  _T_1126; // @[LoadQueue.scala 73:78:@2120.4]
  wire  _T_1127; // @[LoadQueue.scala 73:78:@2121.4]
  wire  _T_1128; // @[LoadQueue.scala 73:78:@2122.4]
  wire  _T_1129; // @[LoadQueue.scala 73:78:@2123.4]
  wire  _T_1130; // @[LoadQueue.scala 73:78:@2124.4]
  wire  _T_1131; // @[LoadQueue.scala 73:78:@2125.4]
  wire  _T_1132; // @[LoadQueue.scala 73:78:@2126.4]
  wire  _T_1133; // @[LoadQueue.scala 73:78:@2127.4]
  wire [2:0] _T_1156; // @[:@2151.6]
  wire [2:0] _GEN_1; // @[LoadQueue.scala 77:20:@2152.6]
  wire [2:0] _GEN_2; // @[LoadQueue.scala 77:20:@2152.6]
  wire [2:0] _GEN_3; // @[LoadQueue.scala 77:20:@2152.6]
  wire [2:0] _GEN_4; // @[LoadQueue.scala 77:20:@2152.6]
  wire [2:0] _GEN_5; // @[LoadQueue.scala 77:20:@2152.6]
  wire [2:0] _GEN_6; // @[LoadQueue.scala 77:20:@2152.6]
  wire [2:0] _GEN_7; // @[LoadQueue.scala 77:20:@2152.6]
  wire [2:0] _GEN_9; // @[LoadQueue.scala 78:18:@2159.6]
  wire [2:0] _GEN_10; // @[LoadQueue.scala 78:18:@2159.6]
  wire [2:0] _GEN_11; // @[LoadQueue.scala 78:18:@2159.6]
  wire [2:0] _GEN_12; // @[LoadQueue.scala 78:18:@2159.6]
  wire [2:0] _GEN_13; // @[LoadQueue.scala 78:18:@2159.6]
  wire [2:0] _GEN_14; // @[LoadQueue.scala 78:18:@2159.6]
  wire [2:0] _GEN_15; // @[LoadQueue.scala 78:18:@2159.6]
  wire [2:0] _GEN_16; // @[LoadQueue.scala 76:25:@2145.4]
  wire [2:0] _GEN_17; // @[LoadQueue.scala 76:25:@2145.4]
  wire [2:0] _T_1174; // @[:@2167.6]
  wire [2:0] _GEN_19; // @[LoadQueue.scala 77:20:@2168.6]
  wire [2:0] _GEN_20; // @[LoadQueue.scala 77:20:@2168.6]
  wire [2:0] _GEN_21; // @[LoadQueue.scala 77:20:@2168.6]
  wire [2:0] _GEN_22; // @[LoadQueue.scala 77:20:@2168.6]
  wire [2:0] _GEN_23; // @[LoadQueue.scala 77:20:@2168.6]
  wire [2:0] _GEN_24; // @[LoadQueue.scala 77:20:@2168.6]
  wire [2:0] _GEN_25; // @[LoadQueue.scala 77:20:@2168.6]
  wire [2:0] _GEN_27; // @[LoadQueue.scala 78:18:@2175.6]
  wire [2:0] _GEN_28; // @[LoadQueue.scala 78:18:@2175.6]
  wire [2:0] _GEN_29; // @[LoadQueue.scala 78:18:@2175.6]
  wire [2:0] _GEN_30; // @[LoadQueue.scala 78:18:@2175.6]
  wire [2:0] _GEN_31; // @[LoadQueue.scala 78:18:@2175.6]
  wire [2:0] _GEN_32; // @[LoadQueue.scala 78:18:@2175.6]
  wire [2:0] _GEN_33; // @[LoadQueue.scala 78:18:@2175.6]
  wire [2:0] _GEN_34; // @[LoadQueue.scala 76:25:@2161.4]
  wire [2:0] _GEN_35; // @[LoadQueue.scala 76:25:@2161.4]
  wire [2:0] _T_1192; // @[:@2183.6]
  wire [2:0] _GEN_37; // @[LoadQueue.scala 77:20:@2184.6]
  wire [2:0] _GEN_38; // @[LoadQueue.scala 77:20:@2184.6]
  wire [2:0] _GEN_39; // @[LoadQueue.scala 77:20:@2184.6]
  wire [2:0] _GEN_40; // @[LoadQueue.scala 77:20:@2184.6]
  wire [2:0] _GEN_41; // @[LoadQueue.scala 77:20:@2184.6]
  wire [2:0] _GEN_42; // @[LoadQueue.scala 77:20:@2184.6]
  wire [2:0] _GEN_43; // @[LoadQueue.scala 77:20:@2184.6]
  wire [2:0] _GEN_45; // @[LoadQueue.scala 78:18:@2191.6]
  wire [2:0] _GEN_46; // @[LoadQueue.scala 78:18:@2191.6]
  wire [2:0] _GEN_47; // @[LoadQueue.scala 78:18:@2191.6]
  wire [2:0] _GEN_48; // @[LoadQueue.scala 78:18:@2191.6]
  wire [2:0] _GEN_49; // @[LoadQueue.scala 78:18:@2191.6]
  wire [2:0] _GEN_50; // @[LoadQueue.scala 78:18:@2191.6]
  wire [2:0] _GEN_51; // @[LoadQueue.scala 78:18:@2191.6]
  wire [2:0] _GEN_52; // @[LoadQueue.scala 76:25:@2177.4]
  wire [2:0] _GEN_53; // @[LoadQueue.scala 76:25:@2177.4]
  wire [2:0] _T_1210; // @[:@2199.6]
  wire [2:0] _GEN_55; // @[LoadQueue.scala 77:20:@2200.6]
  wire [2:0] _GEN_56; // @[LoadQueue.scala 77:20:@2200.6]
  wire [2:0] _GEN_57; // @[LoadQueue.scala 77:20:@2200.6]
  wire [2:0] _GEN_58; // @[LoadQueue.scala 77:20:@2200.6]
  wire [2:0] _GEN_59; // @[LoadQueue.scala 77:20:@2200.6]
  wire [2:0] _GEN_60; // @[LoadQueue.scala 77:20:@2200.6]
  wire [2:0] _GEN_61; // @[LoadQueue.scala 77:20:@2200.6]
  wire [2:0] _GEN_63; // @[LoadQueue.scala 78:18:@2207.6]
  wire [2:0] _GEN_64; // @[LoadQueue.scala 78:18:@2207.6]
  wire [2:0] _GEN_65; // @[LoadQueue.scala 78:18:@2207.6]
  wire [2:0] _GEN_66; // @[LoadQueue.scala 78:18:@2207.6]
  wire [2:0] _GEN_67; // @[LoadQueue.scala 78:18:@2207.6]
  wire [2:0] _GEN_68; // @[LoadQueue.scala 78:18:@2207.6]
  wire [2:0] _GEN_69; // @[LoadQueue.scala 78:18:@2207.6]
  wire [2:0] _GEN_70; // @[LoadQueue.scala 76:25:@2193.4]
  wire [2:0] _GEN_71; // @[LoadQueue.scala 76:25:@2193.4]
  wire [2:0] _T_1228; // @[:@2215.6]
  wire [2:0] _GEN_73; // @[LoadQueue.scala 77:20:@2216.6]
  wire [2:0] _GEN_74; // @[LoadQueue.scala 77:20:@2216.6]
  wire [2:0] _GEN_75; // @[LoadQueue.scala 77:20:@2216.6]
  wire [2:0] _GEN_76; // @[LoadQueue.scala 77:20:@2216.6]
  wire [2:0] _GEN_77; // @[LoadQueue.scala 77:20:@2216.6]
  wire [2:0] _GEN_78; // @[LoadQueue.scala 77:20:@2216.6]
  wire [2:0] _GEN_79; // @[LoadQueue.scala 77:20:@2216.6]
  wire [2:0] _GEN_81; // @[LoadQueue.scala 78:18:@2223.6]
  wire [2:0] _GEN_82; // @[LoadQueue.scala 78:18:@2223.6]
  wire [2:0] _GEN_83; // @[LoadQueue.scala 78:18:@2223.6]
  wire [2:0] _GEN_84; // @[LoadQueue.scala 78:18:@2223.6]
  wire [2:0] _GEN_85; // @[LoadQueue.scala 78:18:@2223.6]
  wire [2:0] _GEN_86; // @[LoadQueue.scala 78:18:@2223.6]
  wire [2:0] _GEN_87; // @[LoadQueue.scala 78:18:@2223.6]
  wire [2:0] _GEN_88; // @[LoadQueue.scala 76:25:@2209.4]
  wire [2:0] _GEN_89; // @[LoadQueue.scala 76:25:@2209.4]
  wire [2:0] _T_1246; // @[:@2231.6]
  wire [2:0] _GEN_91; // @[LoadQueue.scala 77:20:@2232.6]
  wire [2:0] _GEN_92; // @[LoadQueue.scala 77:20:@2232.6]
  wire [2:0] _GEN_93; // @[LoadQueue.scala 77:20:@2232.6]
  wire [2:0] _GEN_94; // @[LoadQueue.scala 77:20:@2232.6]
  wire [2:0] _GEN_95; // @[LoadQueue.scala 77:20:@2232.6]
  wire [2:0] _GEN_96; // @[LoadQueue.scala 77:20:@2232.6]
  wire [2:0] _GEN_97; // @[LoadQueue.scala 77:20:@2232.6]
  wire [2:0] _GEN_99; // @[LoadQueue.scala 78:18:@2239.6]
  wire [2:0] _GEN_100; // @[LoadQueue.scala 78:18:@2239.6]
  wire [2:0] _GEN_101; // @[LoadQueue.scala 78:18:@2239.6]
  wire [2:0] _GEN_102; // @[LoadQueue.scala 78:18:@2239.6]
  wire [2:0] _GEN_103; // @[LoadQueue.scala 78:18:@2239.6]
  wire [2:0] _GEN_104; // @[LoadQueue.scala 78:18:@2239.6]
  wire [2:0] _GEN_105; // @[LoadQueue.scala 78:18:@2239.6]
  wire [2:0] _GEN_106; // @[LoadQueue.scala 76:25:@2225.4]
  wire [2:0] _GEN_107; // @[LoadQueue.scala 76:25:@2225.4]
  wire [2:0] _T_1264; // @[:@2247.6]
  wire [2:0] _GEN_109; // @[LoadQueue.scala 77:20:@2248.6]
  wire [2:0] _GEN_110; // @[LoadQueue.scala 77:20:@2248.6]
  wire [2:0] _GEN_111; // @[LoadQueue.scala 77:20:@2248.6]
  wire [2:0] _GEN_112; // @[LoadQueue.scala 77:20:@2248.6]
  wire [2:0] _GEN_113; // @[LoadQueue.scala 77:20:@2248.6]
  wire [2:0] _GEN_114; // @[LoadQueue.scala 77:20:@2248.6]
  wire [2:0] _GEN_115; // @[LoadQueue.scala 77:20:@2248.6]
  wire [2:0] _GEN_117; // @[LoadQueue.scala 78:18:@2255.6]
  wire [2:0] _GEN_118; // @[LoadQueue.scala 78:18:@2255.6]
  wire [2:0] _GEN_119; // @[LoadQueue.scala 78:18:@2255.6]
  wire [2:0] _GEN_120; // @[LoadQueue.scala 78:18:@2255.6]
  wire [2:0] _GEN_121; // @[LoadQueue.scala 78:18:@2255.6]
  wire [2:0] _GEN_122; // @[LoadQueue.scala 78:18:@2255.6]
  wire [2:0] _GEN_123; // @[LoadQueue.scala 78:18:@2255.6]
  wire [2:0] _GEN_124; // @[LoadQueue.scala 76:25:@2241.4]
  wire [2:0] _GEN_125; // @[LoadQueue.scala 76:25:@2241.4]
  wire [2:0] _T_1282; // @[:@2263.6]
  wire [2:0] _GEN_127; // @[LoadQueue.scala 77:20:@2264.6]
  wire [2:0] _GEN_128; // @[LoadQueue.scala 77:20:@2264.6]
  wire [2:0] _GEN_129; // @[LoadQueue.scala 77:20:@2264.6]
  wire [2:0] _GEN_130; // @[LoadQueue.scala 77:20:@2264.6]
  wire [2:0] _GEN_131; // @[LoadQueue.scala 77:20:@2264.6]
  wire [2:0] _GEN_132; // @[LoadQueue.scala 77:20:@2264.6]
  wire [2:0] _GEN_133; // @[LoadQueue.scala 77:20:@2264.6]
  wire [2:0] _GEN_135; // @[LoadQueue.scala 78:18:@2271.6]
  wire [2:0] _GEN_136; // @[LoadQueue.scala 78:18:@2271.6]
  wire [2:0] _GEN_137; // @[LoadQueue.scala 78:18:@2271.6]
  wire [2:0] _GEN_138; // @[LoadQueue.scala 78:18:@2271.6]
  wire [2:0] _GEN_139; // @[LoadQueue.scala 78:18:@2271.6]
  wire [2:0] _GEN_140; // @[LoadQueue.scala 78:18:@2271.6]
  wire [2:0] _GEN_141; // @[LoadQueue.scala 78:18:@2271.6]
  wire [2:0] _GEN_142; // @[LoadQueue.scala 76:25:@2257.4]
  wire [2:0] _GEN_143; // @[LoadQueue.scala 76:25:@2257.4]
  reg [2:0] previousStoreHead; // @[LoadQueue.scala 93:34:@2273.4]
  reg [31:0] _RAND_82;
  wire [3:0] _T_1304; // @[util.scala 10:8:@2282.6]
  wire [3:0] _GEN_72; // @[util.scala 10:14:@2283.6]
  wire [3:0] _T_1305; // @[util.scala 10:14:@2283.6]
  wire [3:0] _GEN_799; // @[LoadQueue.scala 97:56:@2284.6]
  wire  _T_1306; // @[LoadQueue.scala 97:56:@2284.6]
  wire  _T_1307; // @[LoadQueue.scala 96:50:@2285.6]
  wire  _T_1309; // @[LoadQueue.scala 96:34:@2286.6]
  wire  _T_1311; // @[LoadQueue.scala 101:36:@2294.8]
  wire  _T_1312; // @[LoadQueue.scala 101:86:@2295.8]
  wire  _T_1313; // @[LoadQueue.scala 101:61:@2296.8]
  wire  _T_1315; // @[LoadQueue.scala 103:36:@2301.10]
  wire  _T_1316; // @[LoadQueue.scala 103:69:@2302.10]
  wire  _T_1317; // @[LoadQueue.scala 104:31:@2303.10]
  wire  _T_1318; // @[LoadQueue.scala 103:94:@2304.10]
  wire  _T_1320; // @[LoadQueue.scala 103:54:@2305.10]
  wire  _T_1321; // @[LoadQueue.scala 103:51:@2306.10]
  wire  _GEN_152; // @[LoadQueue.scala 104:53:@2307.10]
  wire  _GEN_153; // @[LoadQueue.scala 101:102:@2297.8]
  wire  _GEN_154; // @[LoadQueue.scala 99:27:@2290.6]
  wire  _GEN_155; // @[LoadQueue.scala 95:34:@2275.4]
  wire [3:0] _T_1334; // @[util.scala 10:8:@2318.6]
  wire [3:0] _GEN_80; // @[util.scala 10:14:@2319.6]
  wire [3:0] _T_1335; // @[util.scala 10:14:@2319.6]
  wire  _T_1336; // @[LoadQueue.scala 97:56:@2320.6]
  wire  _T_1337; // @[LoadQueue.scala 96:50:@2321.6]
  wire  _T_1339; // @[LoadQueue.scala 96:34:@2322.6]
  wire  _T_1341; // @[LoadQueue.scala 101:36:@2330.8]
  wire  _T_1342; // @[LoadQueue.scala 101:86:@2331.8]
  wire  _T_1343; // @[LoadQueue.scala 101:61:@2332.8]
  wire  _T_1346; // @[LoadQueue.scala 103:69:@2338.10]
  wire  _T_1347; // @[LoadQueue.scala 104:31:@2339.10]
  wire  _T_1348; // @[LoadQueue.scala 103:94:@2340.10]
  wire  _T_1350; // @[LoadQueue.scala 103:54:@2341.10]
  wire  _T_1351; // @[LoadQueue.scala 103:51:@2342.10]
  wire  _GEN_164; // @[LoadQueue.scala 104:53:@2343.10]
  wire  _GEN_165; // @[LoadQueue.scala 101:102:@2333.8]
  wire  _GEN_166; // @[LoadQueue.scala 99:27:@2326.6]
  wire  _GEN_167; // @[LoadQueue.scala 95:34:@2311.4]
  wire [3:0] _T_1364; // @[util.scala 10:8:@2354.6]
  wire [3:0] _GEN_90; // @[util.scala 10:14:@2355.6]
  wire [3:0] _T_1365; // @[util.scala 10:14:@2355.6]
  wire  _T_1366; // @[LoadQueue.scala 97:56:@2356.6]
  wire  _T_1367; // @[LoadQueue.scala 96:50:@2357.6]
  wire  _T_1369; // @[LoadQueue.scala 96:34:@2358.6]
  wire  _T_1371; // @[LoadQueue.scala 101:36:@2366.8]
  wire  _T_1372; // @[LoadQueue.scala 101:86:@2367.8]
  wire  _T_1373; // @[LoadQueue.scala 101:61:@2368.8]
  wire  _T_1376; // @[LoadQueue.scala 103:69:@2374.10]
  wire  _T_1377; // @[LoadQueue.scala 104:31:@2375.10]
  wire  _T_1378; // @[LoadQueue.scala 103:94:@2376.10]
  wire  _T_1380; // @[LoadQueue.scala 103:54:@2377.10]
  wire  _T_1381; // @[LoadQueue.scala 103:51:@2378.10]
  wire  _GEN_176; // @[LoadQueue.scala 104:53:@2379.10]
  wire  _GEN_177; // @[LoadQueue.scala 101:102:@2369.8]
  wire  _GEN_178; // @[LoadQueue.scala 99:27:@2362.6]
  wire  _GEN_179; // @[LoadQueue.scala 95:34:@2347.4]
  wire [3:0] _T_1394; // @[util.scala 10:8:@2390.6]
  wire [3:0] _GEN_98; // @[util.scala 10:14:@2391.6]
  wire [3:0] _T_1395; // @[util.scala 10:14:@2391.6]
  wire  _T_1396; // @[LoadQueue.scala 97:56:@2392.6]
  wire  _T_1397; // @[LoadQueue.scala 96:50:@2393.6]
  wire  _T_1399; // @[LoadQueue.scala 96:34:@2394.6]
  wire  _T_1401; // @[LoadQueue.scala 101:36:@2402.8]
  wire  _T_1402; // @[LoadQueue.scala 101:86:@2403.8]
  wire  _T_1403; // @[LoadQueue.scala 101:61:@2404.8]
  wire  _T_1406; // @[LoadQueue.scala 103:69:@2410.10]
  wire  _T_1407; // @[LoadQueue.scala 104:31:@2411.10]
  wire  _T_1408; // @[LoadQueue.scala 103:94:@2412.10]
  wire  _T_1410; // @[LoadQueue.scala 103:54:@2413.10]
  wire  _T_1411; // @[LoadQueue.scala 103:51:@2414.10]
  wire  _GEN_188; // @[LoadQueue.scala 104:53:@2415.10]
  wire  _GEN_189; // @[LoadQueue.scala 101:102:@2405.8]
  wire  _GEN_190; // @[LoadQueue.scala 99:27:@2398.6]
  wire  _GEN_191; // @[LoadQueue.scala 95:34:@2383.4]
  wire [3:0] _T_1424; // @[util.scala 10:8:@2426.6]
  wire [3:0] _GEN_108; // @[util.scala 10:14:@2427.6]
  wire [3:0] _T_1425; // @[util.scala 10:14:@2427.6]
  wire  _T_1426; // @[LoadQueue.scala 97:56:@2428.6]
  wire  _T_1427; // @[LoadQueue.scala 96:50:@2429.6]
  wire  _T_1429; // @[LoadQueue.scala 96:34:@2430.6]
  wire  _T_1431; // @[LoadQueue.scala 101:36:@2438.8]
  wire  _T_1432; // @[LoadQueue.scala 101:86:@2439.8]
  wire  _T_1433; // @[LoadQueue.scala 101:61:@2440.8]
  wire  _T_1436; // @[LoadQueue.scala 103:69:@2446.10]
  wire  _T_1437; // @[LoadQueue.scala 104:31:@2447.10]
  wire  _T_1438; // @[LoadQueue.scala 103:94:@2448.10]
  wire  _T_1440; // @[LoadQueue.scala 103:54:@2449.10]
  wire  _T_1441; // @[LoadQueue.scala 103:51:@2450.10]
  wire  _GEN_200; // @[LoadQueue.scala 104:53:@2451.10]
  wire  _GEN_201; // @[LoadQueue.scala 101:102:@2441.8]
  wire  _GEN_202; // @[LoadQueue.scala 99:27:@2434.6]
  wire  _GEN_203; // @[LoadQueue.scala 95:34:@2419.4]
  wire [3:0] _T_1454; // @[util.scala 10:8:@2462.6]
  wire [3:0] _GEN_116; // @[util.scala 10:14:@2463.6]
  wire [3:0] _T_1455; // @[util.scala 10:14:@2463.6]
  wire  _T_1456; // @[LoadQueue.scala 97:56:@2464.6]
  wire  _T_1457; // @[LoadQueue.scala 96:50:@2465.6]
  wire  _T_1459; // @[LoadQueue.scala 96:34:@2466.6]
  wire  _T_1461; // @[LoadQueue.scala 101:36:@2474.8]
  wire  _T_1462; // @[LoadQueue.scala 101:86:@2475.8]
  wire  _T_1463; // @[LoadQueue.scala 101:61:@2476.8]
  wire  _T_1466; // @[LoadQueue.scala 103:69:@2482.10]
  wire  _T_1467; // @[LoadQueue.scala 104:31:@2483.10]
  wire  _T_1468; // @[LoadQueue.scala 103:94:@2484.10]
  wire  _T_1470; // @[LoadQueue.scala 103:54:@2485.10]
  wire  _T_1471; // @[LoadQueue.scala 103:51:@2486.10]
  wire  _GEN_212; // @[LoadQueue.scala 104:53:@2487.10]
  wire  _GEN_213; // @[LoadQueue.scala 101:102:@2477.8]
  wire  _GEN_214; // @[LoadQueue.scala 99:27:@2470.6]
  wire  _GEN_215; // @[LoadQueue.scala 95:34:@2455.4]
  wire [3:0] _T_1484; // @[util.scala 10:8:@2498.6]
  wire [3:0] _GEN_126; // @[util.scala 10:14:@2499.6]
  wire [3:0] _T_1485; // @[util.scala 10:14:@2499.6]
  wire  _T_1486; // @[LoadQueue.scala 97:56:@2500.6]
  wire  _T_1487; // @[LoadQueue.scala 96:50:@2501.6]
  wire  _T_1489; // @[LoadQueue.scala 96:34:@2502.6]
  wire  _T_1491; // @[LoadQueue.scala 101:36:@2510.8]
  wire  _T_1492; // @[LoadQueue.scala 101:86:@2511.8]
  wire  _T_1493; // @[LoadQueue.scala 101:61:@2512.8]
  wire  _T_1496; // @[LoadQueue.scala 103:69:@2518.10]
  wire  _T_1497; // @[LoadQueue.scala 104:31:@2519.10]
  wire  _T_1498; // @[LoadQueue.scala 103:94:@2520.10]
  wire  _T_1500; // @[LoadQueue.scala 103:54:@2521.10]
  wire  _T_1501; // @[LoadQueue.scala 103:51:@2522.10]
  wire  _GEN_224; // @[LoadQueue.scala 104:53:@2523.10]
  wire  _GEN_225; // @[LoadQueue.scala 101:102:@2513.8]
  wire  _GEN_226; // @[LoadQueue.scala 99:27:@2506.6]
  wire  _GEN_227; // @[LoadQueue.scala 95:34:@2491.4]
  wire [3:0] _T_1514; // @[util.scala 10:8:@2534.6]
  wire [3:0] _GEN_134; // @[util.scala 10:14:@2535.6]
  wire [3:0] _T_1515; // @[util.scala 10:14:@2535.6]
  wire  _T_1516; // @[LoadQueue.scala 97:56:@2536.6]
  wire  _T_1517; // @[LoadQueue.scala 96:50:@2537.6]
  wire  _T_1519; // @[LoadQueue.scala 96:34:@2538.6]
  wire  _T_1521; // @[LoadQueue.scala 101:36:@2546.8]
  wire  _T_1522; // @[LoadQueue.scala 101:86:@2547.8]
  wire  _T_1523; // @[LoadQueue.scala 101:61:@2548.8]
  wire  _T_1526; // @[LoadQueue.scala 103:69:@2554.10]
  wire  _T_1527; // @[LoadQueue.scala 104:31:@2555.10]
  wire  _T_1528; // @[LoadQueue.scala 103:94:@2556.10]
  wire  _T_1530; // @[LoadQueue.scala 103:54:@2557.10]
  wire  _T_1531; // @[LoadQueue.scala 103:51:@2558.10]
  wire  _GEN_236; // @[LoadQueue.scala 104:53:@2559.10]
  wire  _GEN_237; // @[LoadQueue.scala 101:102:@2549.8]
  wire  _GEN_238; // @[LoadQueue.scala 99:27:@2542.6]
  wire  _GEN_239; // @[LoadQueue.scala 95:34:@2527.4]
  wire [7:0] _T_1535; // @[OneHot.scala 52:12:@2564.4]
  wire  _T_1537; // @[util.scala 60:60:@2566.4]
  wire  _T_1538; // @[util.scala 60:60:@2567.4]
  wire  _T_1539; // @[util.scala 60:60:@2568.4]
  wire  _T_1540; // @[util.scala 60:60:@2569.4]
  wire  _T_1541; // @[util.scala 60:60:@2570.4]
  wire  _T_1542; // @[util.scala 60:60:@2571.4]
  wire  _T_1543; // @[util.scala 60:60:@2572.4]
  wire  _T_1544; // @[util.scala 60:60:@2573.4]
  wire [255:0] _T_2323; // @[Mux.scala 19:72:@3025.4]
  wire [255:0] _T_2325; // @[Mux.scala 19:72:@3026.4]
  wire [255:0] _T_2332; // @[Mux.scala 19:72:@3033.4]
  wire [255:0] _T_2334; // @[Mux.scala 19:72:@3034.4]
  wire [255:0] _T_2341; // @[Mux.scala 19:72:@3041.4]
  wire [255:0] _T_2343; // @[Mux.scala 19:72:@3042.4]
  wire [255:0] _T_2350; // @[Mux.scala 19:72:@3049.4]
  wire [255:0] _T_2352; // @[Mux.scala 19:72:@3050.4]
  wire [255:0] _T_2359; // @[Mux.scala 19:72:@3057.4]
  wire [255:0] _T_2361; // @[Mux.scala 19:72:@3058.4]
  wire [255:0] _T_2368; // @[Mux.scala 19:72:@3065.4]
  wire [255:0] _T_2370; // @[Mux.scala 19:72:@3066.4]
  wire [255:0] _T_2377; // @[Mux.scala 19:72:@3073.4]
  wire [255:0] _T_2379; // @[Mux.scala 19:72:@3074.4]
  wire [255:0] _T_2386; // @[Mux.scala 19:72:@3081.4]
  wire [255:0] _T_2388; // @[Mux.scala 19:72:@3082.4]
  wire [255:0] _T_2389; // @[Mux.scala 19:72:@3083.4]
  wire [255:0] _T_2390; // @[Mux.scala 19:72:@3084.4]
  wire [255:0] _T_2391; // @[Mux.scala 19:72:@3085.4]
  wire [255:0] _T_2392; // @[Mux.scala 19:72:@3086.4]
  wire [255:0] _T_2393; // @[Mux.scala 19:72:@3087.4]
  wire [255:0] _T_2394; // @[Mux.scala 19:72:@3088.4]
  wire [255:0] _T_2395; // @[Mux.scala 19:72:@3089.4]
  wire [7:0] _T_2636; // @[Mux.scala 19:72:@3207.4]
  wire [7:0] _T_2638; // @[Mux.scala 19:72:@3208.4]
  wire [7:0] _T_2645; // @[Mux.scala 19:72:@3215.4]
  wire [7:0] _T_2647; // @[Mux.scala 19:72:@3216.4]
  wire [7:0] _T_2654; // @[Mux.scala 19:72:@3223.4]
  wire [7:0] _T_2656; // @[Mux.scala 19:72:@3224.4]
  wire [7:0] _T_2663; // @[Mux.scala 19:72:@3231.4]
  wire [7:0] _T_2665; // @[Mux.scala 19:72:@3232.4]
  wire [7:0] _T_2672; // @[Mux.scala 19:72:@3239.4]
  wire [7:0] _T_2674; // @[Mux.scala 19:72:@3240.4]
  wire [7:0] _T_2681; // @[Mux.scala 19:72:@3247.4]
  wire [7:0] _T_2683; // @[Mux.scala 19:72:@3248.4]
  wire [7:0] _T_2690; // @[Mux.scala 19:72:@3255.4]
  wire [7:0] _T_2692; // @[Mux.scala 19:72:@3256.4]
  wire [7:0] _T_2699; // @[Mux.scala 19:72:@3263.4]
  wire [7:0] _T_2701; // @[Mux.scala 19:72:@3264.4]
  wire [7:0] _T_2702; // @[Mux.scala 19:72:@3265.4]
  wire [7:0] _T_2703; // @[Mux.scala 19:72:@3266.4]
  wire [7:0] _T_2704; // @[Mux.scala 19:72:@3267.4]
  wire [7:0] _T_2705; // @[Mux.scala 19:72:@3268.4]
  wire [7:0] _T_2706; // @[Mux.scala 19:72:@3269.4]
  wire [7:0] _T_2707; // @[Mux.scala 19:72:@3270.4]
  wire [7:0] _T_2708; // @[Mux.scala 19:72:@3271.4]
  wire  _T_2785; // @[LoadQueue.scala 121:105:@3291.4]
  wire  _T_2787; // @[LoadQueue.scala 122:18:@3292.4]
  wire  _T_2789; // @[LoadQueue.scala 122:36:@3293.4]
  wire  _T_2790; // @[LoadQueue.scala 122:27:@3294.4]
  wire  _T_2792; // @[LoadQueue.scala 122:52:@3295.4]
  wire  _T_2794; // @[LoadQueue.scala 122:85:@3296.4]
  wire  _T_2796; // @[LoadQueue.scala 122:103:@3297.4]
  wire  _T_2797; // @[LoadQueue.scala 122:94:@3298.4]
  wire  _T_2799; // @[LoadQueue.scala 122:70:@3299.4]
  wire  _T_2800; // @[LoadQueue.scala 122:67:@3300.4]
  wire  validEntriesInStoreQ_0; // @[LoadQueue.scala 121:91:@3301.4]
  wire  _T_2804; // @[LoadQueue.scala 122:18:@3303.4]
  wire  _T_2806; // @[LoadQueue.scala 122:36:@3304.4]
  wire  _T_2807; // @[LoadQueue.scala 122:27:@3305.4]
  wire  _T_2811; // @[LoadQueue.scala 122:85:@3307.4]
  wire  _T_2813; // @[LoadQueue.scala 122:103:@3308.4]
  wire  _T_2814; // @[LoadQueue.scala 122:94:@3309.4]
  wire  _T_2816; // @[LoadQueue.scala 122:70:@3310.4]
  wire  _T_2817; // @[LoadQueue.scala 122:67:@3311.4]
  wire  validEntriesInStoreQ_1; // @[LoadQueue.scala 121:91:@3312.4]
  wire  _T_2821; // @[LoadQueue.scala 122:18:@3314.4]
  wire  _T_2823; // @[LoadQueue.scala 122:36:@3315.4]
  wire  _T_2824; // @[LoadQueue.scala 122:27:@3316.4]
  wire  _T_2828; // @[LoadQueue.scala 122:85:@3318.4]
  wire  _T_2830; // @[LoadQueue.scala 122:103:@3319.4]
  wire  _T_2831; // @[LoadQueue.scala 122:94:@3320.4]
  wire  _T_2833; // @[LoadQueue.scala 122:70:@3321.4]
  wire  _T_2834; // @[LoadQueue.scala 122:67:@3322.4]
  wire  validEntriesInStoreQ_2; // @[LoadQueue.scala 121:91:@3323.4]
  wire  _T_2838; // @[LoadQueue.scala 122:18:@3325.4]
  wire  _T_2840; // @[LoadQueue.scala 122:36:@3326.4]
  wire  _T_2841; // @[LoadQueue.scala 122:27:@3327.4]
  wire  _T_2845; // @[LoadQueue.scala 122:85:@3329.4]
  wire  _T_2847; // @[LoadQueue.scala 122:103:@3330.4]
  wire  _T_2848; // @[LoadQueue.scala 122:94:@3331.4]
  wire  _T_2850; // @[LoadQueue.scala 122:70:@3332.4]
  wire  _T_2851; // @[LoadQueue.scala 122:67:@3333.4]
  wire  validEntriesInStoreQ_3; // @[LoadQueue.scala 121:91:@3334.4]
  wire  _T_2855; // @[LoadQueue.scala 122:18:@3336.4]
  wire  _T_2857; // @[LoadQueue.scala 122:36:@3337.4]
  wire  _T_2858; // @[LoadQueue.scala 122:27:@3338.4]
  wire  _T_2862; // @[LoadQueue.scala 122:85:@3340.4]
  wire  _T_2864; // @[LoadQueue.scala 122:103:@3341.4]
  wire  _T_2865; // @[LoadQueue.scala 122:94:@3342.4]
  wire  _T_2867; // @[LoadQueue.scala 122:70:@3343.4]
  wire  _T_2868; // @[LoadQueue.scala 122:67:@3344.4]
  wire  validEntriesInStoreQ_4; // @[LoadQueue.scala 121:91:@3345.4]
  wire  _T_2872; // @[LoadQueue.scala 122:18:@3347.4]
  wire  _T_2874; // @[LoadQueue.scala 122:36:@3348.4]
  wire  _T_2875; // @[LoadQueue.scala 122:27:@3349.4]
  wire  _T_2879; // @[LoadQueue.scala 122:85:@3351.4]
  wire  _T_2881; // @[LoadQueue.scala 122:103:@3352.4]
  wire  _T_2882; // @[LoadQueue.scala 122:94:@3353.4]
  wire  _T_2884; // @[LoadQueue.scala 122:70:@3354.4]
  wire  _T_2885; // @[LoadQueue.scala 122:67:@3355.4]
  wire  validEntriesInStoreQ_5; // @[LoadQueue.scala 121:91:@3356.4]
  wire  _T_2889; // @[LoadQueue.scala 122:18:@3358.4]
  wire  _T_2891; // @[LoadQueue.scala 122:36:@3359.4]
  wire  _T_2892; // @[LoadQueue.scala 122:27:@3360.4]
  wire  _T_2896; // @[LoadQueue.scala 122:85:@3362.4]
  wire  _T_2898; // @[LoadQueue.scala 122:103:@3363.4]
  wire  _T_2899; // @[LoadQueue.scala 122:94:@3364.4]
  wire  _T_2901; // @[LoadQueue.scala 122:70:@3365.4]
  wire  _T_2902; // @[LoadQueue.scala 122:67:@3366.4]
  wire  validEntriesInStoreQ_6; // @[LoadQueue.scala 121:91:@3367.4]
  wire  validEntriesInStoreQ_7; // @[LoadQueue.scala 121:91:@3378.4]
  wire  storesToCheck_0_0; // @[LoadQueue.scala 131:10:@3397.4]
  wire  _T_3318; // @[LoadQueue.scala 131:81:@3400.4]
  wire  _T_3319; // @[LoadQueue.scala 131:72:@3401.4]
  wire  _T_3321; // @[LoadQueue.scala 132:33:@3402.4]
  wire  _T_3324; // @[LoadQueue.scala 132:41:@3404.4]
  wire  _T_3326; // @[LoadQueue.scala 132:9:@3405.4]
  wire  storesToCheck_0_1; // @[LoadQueue.scala 131:10:@3406.4]
  wire  _T_3332; // @[LoadQueue.scala 131:81:@3409.4]
  wire  _T_3333; // @[LoadQueue.scala 131:72:@3410.4]
  wire  _T_3335; // @[LoadQueue.scala 132:33:@3411.4]
  wire  _T_3338; // @[LoadQueue.scala 132:41:@3413.4]
  wire  _T_3340; // @[LoadQueue.scala 132:9:@3414.4]
  wire  storesToCheck_0_2; // @[LoadQueue.scala 131:10:@3415.4]
  wire  _T_3346; // @[LoadQueue.scala 131:81:@3418.4]
  wire  _T_3347; // @[LoadQueue.scala 131:72:@3419.4]
  wire  _T_3349; // @[LoadQueue.scala 132:33:@3420.4]
  wire  _T_3352; // @[LoadQueue.scala 132:41:@3422.4]
  wire  _T_3354; // @[LoadQueue.scala 132:9:@3423.4]
  wire  storesToCheck_0_3; // @[LoadQueue.scala 131:10:@3424.4]
  wire  _T_3360; // @[LoadQueue.scala 131:81:@3427.4]
  wire  _T_3361; // @[LoadQueue.scala 131:72:@3428.4]
  wire  _T_3363; // @[LoadQueue.scala 132:33:@3429.4]
  wire  _T_3366; // @[LoadQueue.scala 132:41:@3431.4]
  wire  _T_3368; // @[LoadQueue.scala 132:9:@3432.4]
  wire  storesToCheck_0_4; // @[LoadQueue.scala 131:10:@3433.4]
  wire  _T_3374; // @[LoadQueue.scala 131:81:@3436.4]
  wire  _T_3375; // @[LoadQueue.scala 131:72:@3437.4]
  wire  _T_3377; // @[LoadQueue.scala 132:33:@3438.4]
  wire  _T_3380; // @[LoadQueue.scala 132:41:@3440.4]
  wire  _T_3382; // @[LoadQueue.scala 132:9:@3441.4]
  wire  storesToCheck_0_5; // @[LoadQueue.scala 131:10:@3442.4]
  wire  _T_3388; // @[LoadQueue.scala 131:81:@3445.4]
  wire  _T_3389; // @[LoadQueue.scala 131:72:@3446.4]
  wire  _T_3391; // @[LoadQueue.scala 132:33:@3447.4]
  wire  _T_3394; // @[LoadQueue.scala 132:41:@3449.4]
  wire  _T_3396; // @[LoadQueue.scala 132:9:@3450.4]
  wire  storesToCheck_0_6; // @[LoadQueue.scala 131:10:@3451.4]
  wire  _T_3402; // @[LoadQueue.scala 131:81:@3454.4]
  wire  storesToCheck_0_7; // @[LoadQueue.scala 131:10:@3460.4]
  wire  storesToCheck_1_0; // @[LoadQueue.scala 131:10:@3486.4]
  wire  _T_3444; // @[LoadQueue.scala 131:81:@3489.4]
  wire  _T_3445; // @[LoadQueue.scala 131:72:@3490.4]
  wire  _T_3447; // @[LoadQueue.scala 132:33:@3491.4]
  wire  _T_3450; // @[LoadQueue.scala 132:41:@3493.4]
  wire  _T_3452; // @[LoadQueue.scala 132:9:@3494.4]
  wire  storesToCheck_1_1; // @[LoadQueue.scala 131:10:@3495.4]
  wire  _T_3458; // @[LoadQueue.scala 131:81:@3498.4]
  wire  _T_3459; // @[LoadQueue.scala 131:72:@3499.4]
  wire  _T_3461; // @[LoadQueue.scala 132:33:@3500.4]
  wire  _T_3464; // @[LoadQueue.scala 132:41:@3502.4]
  wire  _T_3466; // @[LoadQueue.scala 132:9:@3503.4]
  wire  storesToCheck_1_2; // @[LoadQueue.scala 131:10:@3504.4]
  wire  _T_3472; // @[LoadQueue.scala 131:81:@3507.4]
  wire  _T_3473; // @[LoadQueue.scala 131:72:@3508.4]
  wire  _T_3475; // @[LoadQueue.scala 132:33:@3509.4]
  wire  _T_3478; // @[LoadQueue.scala 132:41:@3511.4]
  wire  _T_3480; // @[LoadQueue.scala 132:9:@3512.4]
  wire  storesToCheck_1_3; // @[LoadQueue.scala 131:10:@3513.4]
  wire  _T_3486; // @[LoadQueue.scala 131:81:@3516.4]
  wire  _T_3487; // @[LoadQueue.scala 131:72:@3517.4]
  wire  _T_3489; // @[LoadQueue.scala 132:33:@3518.4]
  wire  _T_3492; // @[LoadQueue.scala 132:41:@3520.4]
  wire  _T_3494; // @[LoadQueue.scala 132:9:@3521.4]
  wire  storesToCheck_1_4; // @[LoadQueue.scala 131:10:@3522.4]
  wire  _T_3500; // @[LoadQueue.scala 131:81:@3525.4]
  wire  _T_3501; // @[LoadQueue.scala 131:72:@3526.4]
  wire  _T_3503; // @[LoadQueue.scala 132:33:@3527.4]
  wire  _T_3506; // @[LoadQueue.scala 132:41:@3529.4]
  wire  _T_3508; // @[LoadQueue.scala 132:9:@3530.4]
  wire  storesToCheck_1_5; // @[LoadQueue.scala 131:10:@3531.4]
  wire  _T_3514; // @[LoadQueue.scala 131:81:@3534.4]
  wire  _T_3515; // @[LoadQueue.scala 131:72:@3535.4]
  wire  _T_3517; // @[LoadQueue.scala 132:33:@3536.4]
  wire  _T_3520; // @[LoadQueue.scala 132:41:@3538.4]
  wire  _T_3522; // @[LoadQueue.scala 132:9:@3539.4]
  wire  storesToCheck_1_6; // @[LoadQueue.scala 131:10:@3540.4]
  wire  _T_3528; // @[LoadQueue.scala 131:81:@3543.4]
  wire  storesToCheck_1_7; // @[LoadQueue.scala 131:10:@3549.4]
  wire  storesToCheck_2_0; // @[LoadQueue.scala 131:10:@3575.4]
  wire  _T_3570; // @[LoadQueue.scala 131:81:@3578.4]
  wire  _T_3571; // @[LoadQueue.scala 131:72:@3579.4]
  wire  _T_3573; // @[LoadQueue.scala 132:33:@3580.4]
  wire  _T_3576; // @[LoadQueue.scala 132:41:@3582.4]
  wire  _T_3578; // @[LoadQueue.scala 132:9:@3583.4]
  wire  storesToCheck_2_1; // @[LoadQueue.scala 131:10:@3584.4]
  wire  _T_3584; // @[LoadQueue.scala 131:81:@3587.4]
  wire  _T_3585; // @[LoadQueue.scala 131:72:@3588.4]
  wire  _T_3587; // @[LoadQueue.scala 132:33:@3589.4]
  wire  _T_3590; // @[LoadQueue.scala 132:41:@3591.4]
  wire  _T_3592; // @[LoadQueue.scala 132:9:@3592.4]
  wire  storesToCheck_2_2; // @[LoadQueue.scala 131:10:@3593.4]
  wire  _T_3598; // @[LoadQueue.scala 131:81:@3596.4]
  wire  _T_3599; // @[LoadQueue.scala 131:72:@3597.4]
  wire  _T_3601; // @[LoadQueue.scala 132:33:@3598.4]
  wire  _T_3604; // @[LoadQueue.scala 132:41:@3600.4]
  wire  _T_3606; // @[LoadQueue.scala 132:9:@3601.4]
  wire  storesToCheck_2_3; // @[LoadQueue.scala 131:10:@3602.4]
  wire  _T_3612; // @[LoadQueue.scala 131:81:@3605.4]
  wire  _T_3613; // @[LoadQueue.scala 131:72:@3606.4]
  wire  _T_3615; // @[LoadQueue.scala 132:33:@3607.4]
  wire  _T_3618; // @[LoadQueue.scala 132:41:@3609.4]
  wire  _T_3620; // @[LoadQueue.scala 132:9:@3610.4]
  wire  storesToCheck_2_4; // @[LoadQueue.scala 131:10:@3611.4]
  wire  _T_3626; // @[LoadQueue.scala 131:81:@3614.4]
  wire  _T_3627; // @[LoadQueue.scala 131:72:@3615.4]
  wire  _T_3629; // @[LoadQueue.scala 132:33:@3616.4]
  wire  _T_3632; // @[LoadQueue.scala 132:41:@3618.4]
  wire  _T_3634; // @[LoadQueue.scala 132:9:@3619.4]
  wire  storesToCheck_2_5; // @[LoadQueue.scala 131:10:@3620.4]
  wire  _T_3640; // @[LoadQueue.scala 131:81:@3623.4]
  wire  _T_3641; // @[LoadQueue.scala 131:72:@3624.4]
  wire  _T_3643; // @[LoadQueue.scala 132:33:@3625.4]
  wire  _T_3646; // @[LoadQueue.scala 132:41:@3627.4]
  wire  _T_3648; // @[LoadQueue.scala 132:9:@3628.4]
  wire  storesToCheck_2_6; // @[LoadQueue.scala 131:10:@3629.4]
  wire  _T_3654; // @[LoadQueue.scala 131:81:@3632.4]
  wire  storesToCheck_2_7; // @[LoadQueue.scala 131:10:@3638.4]
  wire  storesToCheck_3_0; // @[LoadQueue.scala 131:10:@3664.4]
  wire  _T_3696; // @[LoadQueue.scala 131:81:@3667.4]
  wire  _T_3697; // @[LoadQueue.scala 131:72:@3668.4]
  wire  _T_3699; // @[LoadQueue.scala 132:33:@3669.4]
  wire  _T_3702; // @[LoadQueue.scala 132:41:@3671.4]
  wire  _T_3704; // @[LoadQueue.scala 132:9:@3672.4]
  wire  storesToCheck_3_1; // @[LoadQueue.scala 131:10:@3673.4]
  wire  _T_3710; // @[LoadQueue.scala 131:81:@3676.4]
  wire  _T_3711; // @[LoadQueue.scala 131:72:@3677.4]
  wire  _T_3713; // @[LoadQueue.scala 132:33:@3678.4]
  wire  _T_3716; // @[LoadQueue.scala 132:41:@3680.4]
  wire  _T_3718; // @[LoadQueue.scala 132:9:@3681.4]
  wire  storesToCheck_3_2; // @[LoadQueue.scala 131:10:@3682.4]
  wire  _T_3724; // @[LoadQueue.scala 131:81:@3685.4]
  wire  _T_3725; // @[LoadQueue.scala 131:72:@3686.4]
  wire  _T_3727; // @[LoadQueue.scala 132:33:@3687.4]
  wire  _T_3730; // @[LoadQueue.scala 132:41:@3689.4]
  wire  _T_3732; // @[LoadQueue.scala 132:9:@3690.4]
  wire  storesToCheck_3_3; // @[LoadQueue.scala 131:10:@3691.4]
  wire  _T_3738; // @[LoadQueue.scala 131:81:@3694.4]
  wire  _T_3739; // @[LoadQueue.scala 131:72:@3695.4]
  wire  _T_3741; // @[LoadQueue.scala 132:33:@3696.4]
  wire  _T_3744; // @[LoadQueue.scala 132:41:@3698.4]
  wire  _T_3746; // @[LoadQueue.scala 132:9:@3699.4]
  wire  storesToCheck_3_4; // @[LoadQueue.scala 131:10:@3700.4]
  wire  _T_3752; // @[LoadQueue.scala 131:81:@3703.4]
  wire  _T_3753; // @[LoadQueue.scala 131:72:@3704.4]
  wire  _T_3755; // @[LoadQueue.scala 132:33:@3705.4]
  wire  _T_3758; // @[LoadQueue.scala 132:41:@3707.4]
  wire  _T_3760; // @[LoadQueue.scala 132:9:@3708.4]
  wire  storesToCheck_3_5; // @[LoadQueue.scala 131:10:@3709.4]
  wire  _T_3766; // @[LoadQueue.scala 131:81:@3712.4]
  wire  _T_3767; // @[LoadQueue.scala 131:72:@3713.4]
  wire  _T_3769; // @[LoadQueue.scala 132:33:@3714.4]
  wire  _T_3772; // @[LoadQueue.scala 132:41:@3716.4]
  wire  _T_3774; // @[LoadQueue.scala 132:9:@3717.4]
  wire  storesToCheck_3_6; // @[LoadQueue.scala 131:10:@3718.4]
  wire  _T_3780; // @[LoadQueue.scala 131:81:@3721.4]
  wire  storesToCheck_3_7; // @[LoadQueue.scala 131:10:@3727.4]
  wire  storesToCheck_4_0; // @[LoadQueue.scala 131:10:@3753.4]
  wire  _T_3822; // @[LoadQueue.scala 131:81:@3756.4]
  wire  _T_3823; // @[LoadQueue.scala 131:72:@3757.4]
  wire  _T_3825; // @[LoadQueue.scala 132:33:@3758.4]
  wire  _T_3828; // @[LoadQueue.scala 132:41:@3760.4]
  wire  _T_3830; // @[LoadQueue.scala 132:9:@3761.4]
  wire  storesToCheck_4_1; // @[LoadQueue.scala 131:10:@3762.4]
  wire  _T_3836; // @[LoadQueue.scala 131:81:@3765.4]
  wire  _T_3837; // @[LoadQueue.scala 131:72:@3766.4]
  wire  _T_3839; // @[LoadQueue.scala 132:33:@3767.4]
  wire  _T_3842; // @[LoadQueue.scala 132:41:@3769.4]
  wire  _T_3844; // @[LoadQueue.scala 132:9:@3770.4]
  wire  storesToCheck_4_2; // @[LoadQueue.scala 131:10:@3771.4]
  wire  _T_3850; // @[LoadQueue.scala 131:81:@3774.4]
  wire  _T_3851; // @[LoadQueue.scala 131:72:@3775.4]
  wire  _T_3853; // @[LoadQueue.scala 132:33:@3776.4]
  wire  _T_3856; // @[LoadQueue.scala 132:41:@3778.4]
  wire  _T_3858; // @[LoadQueue.scala 132:9:@3779.4]
  wire  storesToCheck_4_3; // @[LoadQueue.scala 131:10:@3780.4]
  wire  _T_3864; // @[LoadQueue.scala 131:81:@3783.4]
  wire  _T_3865; // @[LoadQueue.scala 131:72:@3784.4]
  wire  _T_3867; // @[LoadQueue.scala 132:33:@3785.4]
  wire  _T_3870; // @[LoadQueue.scala 132:41:@3787.4]
  wire  _T_3872; // @[LoadQueue.scala 132:9:@3788.4]
  wire  storesToCheck_4_4; // @[LoadQueue.scala 131:10:@3789.4]
  wire  _T_3878; // @[LoadQueue.scala 131:81:@3792.4]
  wire  _T_3879; // @[LoadQueue.scala 131:72:@3793.4]
  wire  _T_3881; // @[LoadQueue.scala 132:33:@3794.4]
  wire  _T_3884; // @[LoadQueue.scala 132:41:@3796.4]
  wire  _T_3886; // @[LoadQueue.scala 132:9:@3797.4]
  wire  storesToCheck_4_5; // @[LoadQueue.scala 131:10:@3798.4]
  wire  _T_3892; // @[LoadQueue.scala 131:81:@3801.4]
  wire  _T_3893; // @[LoadQueue.scala 131:72:@3802.4]
  wire  _T_3895; // @[LoadQueue.scala 132:33:@3803.4]
  wire  _T_3898; // @[LoadQueue.scala 132:41:@3805.4]
  wire  _T_3900; // @[LoadQueue.scala 132:9:@3806.4]
  wire  storesToCheck_4_6; // @[LoadQueue.scala 131:10:@3807.4]
  wire  _T_3906; // @[LoadQueue.scala 131:81:@3810.4]
  wire  storesToCheck_4_7; // @[LoadQueue.scala 131:10:@3816.4]
  wire  storesToCheck_5_0; // @[LoadQueue.scala 131:10:@3842.4]
  wire  _T_3948; // @[LoadQueue.scala 131:81:@3845.4]
  wire  _T_3949; // @[LoadQueue.scala 131:72:@3846.4]
  wire  _T_3951; // @[LoadQueue.scala 132:33:@3847.4]
  wire  _T_3954; // @[LoadQueue.scala 132:41:@3849.4]
  wire  _T_3956; // @[LoadQueue.scala 132:9:@3850.4]
  wire  storesToCheck_5_1; // @[LoadQueue.scala 131:10:@3851.4]
  wire  _T_3962; // @[LoadQueue.scala 131:81:@3854.4]
  wire  _T_3963; // @[LoadQueue.scala 131:72:@3855.4]
  wire  _T_3965; // @[LoadQueue.scala 132:33:@3856.4]
  wire  _T_3968; // @[LoadQueue.scala 132:41:@3858.4]
  wire  _T_3970; // @[LoadQueue.scala 132:9:@3859.4]
  wire  storesToCheck_5_2; // @[LoadQueue.scala 131:10:@3860.4]
  wire  _T_3976; // @[LoadQueue.scala 131:81:@3863.4]
  wire  _T_3977; // @[LoadQueue.scala 131:72:@3864.4]
  wire  _T_3979; // @[LoadQueue.scala 132:33:@3865.4]
  wire  _T_3982; // @[LoadQueue.scala 132:41:@3867.4]
  wire  _T_3984; // @[LoadQueue.scala 132:9:@3868.4]
  wire  storesToCheck_5_3; // @[LoadQueue.scala 131:10:@3869.4]
  wire  _T_3990; // @[LoadQueue.scala 131:81:@3872.4]
  wire  _T_3991; // @[LoadQueue.scala 131:72:@3873.4]
  wire  _T_3993; // @[LoadQueue.scala 132:33:@3874.4]
  wire  _T_3996; // @[LoadQueue.scala 132:41:@3876.4]
  wire  _T_3998; // @[LoadQueue.scala 132:9:@3877.4]
  wire  storesToCheck_5_4; // @[LoadQueue.scala 131:10:@3878.4]
  wire  _T_4004; // @[LoadQueue.scala 131:81:@3881.4]
  wire  _T_4005; // @[LoadQueue.scala 131:72:@3882.4]
  wire  _T_4007; // @[LoadQueue.scala 132:33:@3883.4]
  wire  _T_4010; // @[LoadQueue.scala 132:41:@3885.4]
  wire  _T_4012; // @[LoadQueue.scala 132:9:@3886.4]
  wire  storesToCheck_5_5; // @[LoadQueue.scala 131:10:@3887.4]
  wire  _T_4018; // @[LoadQueue.scala 131:81:@3890.4]
  wire  _T_4019; // @[LoadQueue.scala 131:72:@3891.4]
  wire  _T_4021; // @[LoadQueue.scala 132:33:@3892.4]
  wire  _T_4024; // @[LoadQueue.scala 132:41:@3894.4]
  wire  _T_4026; // @[LoadQueue.scala 132:9:@3895.4]
  wire  storesToCheck_5_6; // @[LoadQueue.scala 131:10:@3896.4]
  wire  _T_4032; // @[LoadQueue.scala 131:81:@3899.4]
  wire  storesToCheck_5_7; // @[LoadQueue.scala 131:10:@3905.4]
  wire  storesToCheck_6_0; // @[LoadQueue.scala 131:10:@3931.4]
  wire  _T_4074; // @[LoadQueue.scala 131:81:@3934.4]
  wire  _T_4075; // @[LoadQueue.scala 131:72:@3935.4]
  wire  _T_4077; // @[LoadQueue.scala 132:33:@3936.4]
  wire  _T_4080; // @[LoadQueue.scala 132:41:@3938.4]
  wire  _T_4082; // @[LoadQueue.scala 132:9:@3939.4]
  wire  storesToCheck_6_1; // @[LoadQueue.scala 131:10:@3940.4]
  wire  _T_4088; // @[LoadQueue.scala 131:81:@3943.4]
  wire  _T_4089; // @[LoadQueue.scala 131:72:@3944.4]
  wire  _T_4091; // @[LoadQueue.scala 132:33:@3945.4]
  wire  _T_4094; // @[LoadQueue.scala 132:41:@3947.4]
  wire  _T_4096; // @[LoadQueue.scala 132:9:@3948.4]
  wire  storesToCheck_6_2; // @[LoadQueue.scala 131:10:@3949.4]
  wire  _T_4102; // @[LoadQueue.scala 131:81:@3952.4]
  wire  _T_4103; // @[LoadQueue.scala 131:72:@3953.4]
  wire  _T_4105; // @[LoadQueue.scala 132:33:@3954.4]
  wire  _T_4108; // @[LoadQueue.scala 132:41:@3956.4]
  wire  _T_4110; // @[LoadQueue.scala 132:9:@3957.4]
  wire  storesToCheck_6_3; // @[LoadQueue.scala 131:10:@3958.4]
  wire  _T_4116; // @[LoadQueue.scala 131:81:@3961.4]
  wire  _T_4117; // @[LoadQueue.scala 131:72:@3962.4]
  wire  _T_4119; // @[LoadQueue.scala 132:33:@3963.4]
  wire  _T_4122; // @[LoadQueue.scala 132:41:@3965.4]
  wire  _T_4124; // @[LoadQueue.scala 132:9:@3966.4]
  wire  storesToCheck_6_4; // @[LoadQueue.scala 131:10:@3967.4]
  wire  _T_4130; // @[LoadQueue.scala 131:81:@3970.4]
  wire  _T_4131; // @[LoadQueue.scala 131:72:@3971.4]
  wire  _T_4133; // @[LoadQueue.scala 132:33:@3972.4]
  wire  _T_4136; // @[LoadQueue.scala 132:41:@3974.4]
  wire  _T_4138; // @[LoadQueue.scala 132:9:@3975.4]
  wire  storesToCheck_6_5; // @[LoadQueue.scala 131:10:@3976.4]
  wire  _T_4144; // @[LoadQueue.scala 131:81:@3979.4]
  wire  _T_4145; // @[LoadQueue.scala 131:72:@3980.4]
  wire  _T_4147; // @[LoadQueue.scala 132:33:@3981.4]
  wire  _T_4150; // @[LoadQueue.scala 132:41:@3983.4]
  wire  _T_4152; // @[LoadQueue.scala 132:9:@3984.4]
  wire  storesToCheck_6_6; // @[LoadQueue.scala 131:10:@3985.4]
  wire  _T_4158; // @[LoadQueue.scala 131:81:@3988.4]
  wire  storesToCheck_6_7; // @[LoadQueue.scala 131:10:@3994.4]
  wire  storesToCheck_7_0; // @[LoadQueue.scala 131:10:@4020.4]
  wire  _T_4200; // @[LoadQueue.scala 131:81:@4023.4]
  wire  _T_4201; // @[LoadQueue.scala 131:72:@4024.4]
  wire  _T_4203; // @[LoadQueue.scala 132:33:@4025.4]
  wire  _T_4206; // @[LoadQueue.scala 132:41:@4027.4]
  wire  _T_4208; // @[LoadQueue.scala 132:9:@4028.4]
  wire  storesToCheck_7_1; // @[LoadQueue.scala 131:10:@4029.4]
  wire  _T_4214; // @[LoadQueue.scala 131:81:@4032.4]
  wire  _T_4215; // @[LoadQueue.scala 131:72:@4033.4]
  wire  _T_4217; // @[LoadQueue.scala 132:33:@4034.4]
  wire  _T_4220; // @[LoadQueue.scala 132:41:@4036.4]
  wire  _T_4222; // @[LoadQueue.scala 132:9:@4037.4]
  wire  storesToCheck_7_2; // @[LoadQueue.scala 131:10:@4038.4]
  wire  _T_4228; // @[LoadQueue.scala 131:81:@4041.4]
  wire  _T_4229; // @[LoadQueue.scala 131:72:@4042.4]
  wire  _T_4231; // @[LoadQueue.scala 132:33:@4043.4]
  wire  _T_4234; // @[LoadQueue.scala 132:41:@4045.4]
  wire  _T_4236; // @[LoadQueue.scala 132:9:@4046.4]
  wire  storesToCheck_7_3; // @[LoadQueue.scala 131:10:@4047.4]
  wire  _T_4242; // @[LoadQueue.scala 131:81:@4050.4]
  wire  _T_4243; // @[LoadQueue.scala 131:72:@4051.4]
  wire  _T_4245; // @[LoadQueue.scala 132:33:@4052.4]
  wire  _T_4248; // @[LoadQueue.scala 132:41:@4054.4]
  wire  _T_4250; // @[LoadQueue.scala 132:9:@4055.4]
  wire  storesToCheck_7_4; // @[LoadQueue.scala 131:10:@4056.4]
  wire  _T_4256; // @[LoadQueue.scala 131:81:@4059.4]
  wire  _T_4257; // @[LoadQueue.scala 131:72:@4060.4]
  wire  _T_4259; // @[LoadQueue.scala 132:33:@4061.4]
  wire  _T_4262; // @[LoadQueue.scala 132:41:@4063.4]
  wire  _T_4264; // @[LoadQueue.scala 132:9:@4064.4]
  wire  storesToCheck_7_5; // @[LoadQueue.scala 131:10:@4065.4]
  wire  _T_4270; // @[LoadQueue.scala 131:81:@4068.4]
  wire  _T_4271; // @[LoadQueue.scala 131:72:@4069.4]
  wire  _T_4273; // @[LoadQueue.scala 132:33:@4070.4]
  wire  _T_4276; // @[LoadQueue.scala 132:41:@4072.4]
  wire  _T_4278; // @[LoadQueue.scala 132:9:@4073.4]
  wire  storesToCheck_7_6; // @[LoadQueue.scala 131:10:@4074.4]
  wire  _T_4284; // @[LoadQueue.scala 131:81:@4077.4]
  wire  storesToCheck_7_7; // @[LoadQueue.scala 131:10:@4083.4]
  wire  _T_4674; // @[LoadQueue.scala 141:18:@4102.4]
  wire  entriesToCheck_0_0; // @[LoadQueue.scala 141:26:@4103.4]
  wire  _T_4676; // @[LoadQueue.scala 141:18:@4104.4]
  wire  entriesToCheck_0_1; // @[LoadQueue.scala 141:26:@4105.4]
  wire  _T_4678; // @[LoadQueue.scala 141:18:@4106.4]
  wire  entriesToCheck_0_2; // @[LoadQueue.scala 141:26:@4107.4]
  wire  _T_4680; // @[LoadQueue.scala 141:18:@4108.4]
  wire  entriesToCheck_0_3; // @[LoadQueue.scala 141:26:@4109.4]
  wire  _T_4682; // @[LoadQueue.scala 141:18:@4110.4]
  wire  entriesToCheck_0_4; // @[LoadQueue.scala 141:26:@4111.4]
  wire  _T_4684; // @[LoadQueue.scala 141:18:@4112.4]
  wire  entriesToCheck_0_5; // @[LoadQueue.scala 141:26:@4113.4]
  wire  _T_4686; // @[LoadQueue.scala 141:18:@4114.4]
  wire  entriesToCheck_0_6; // @[LoadQueue.scala 141:26:@4115.4]
  wire  _T_4688; // @[LoadQueue.scala 141:18:@4116.4]
  wire  entriesToCheck_0_7; // @[LoadQueue.scala 141:26:@4117.4]
  wire  _T_4690; // @[LoadQueue.scala 141:18:@4126.4]
  wire  entriesToCheck_1_0; // @[LoadQueue.scala 141:26:@4127.4]
  wire  _T_4692; // @[LoadQueue.scala 141:18:@4128.4]
  wire  entriesToCheck_1_1; // @[LoadQueue.scala 141:26:@4129.4]
  wire  _T_4694; // @[LoadQueue.scala 141:18:@4130.4]
  wire  entriesToCheck_1_2; // @[LoadQueue.scala 141:26:@4131.4]
  wire  _T_4696; // @[LoadQueue.scala 141:18:@4132.4]
  wire  entriesToCheck_1_3; // @[LoadQueue.scala 141:26:@4133.4]
  wire  _T_4698; // @[LoadQueue.scala 141:18:@4134.4]
  wire  entriesToCheck_1_4; // @[LoadQueue.scala 141:26:@4135.4]
  wire  _T_4700; // @[LoadQueue.scala 141:18:@4136.4]
  wire  entriesToCheck_1_5; // @[LoadQueue.scala 141:26:@4137.4]
  wire  _T_4702; // @[LoadQueue.scala 141:18:@4138.4]
  wire  entriesToCheck_1_6; // @[LoadQueue.scala 141:26:@4139.4]
  wire  _T_4704; // @[LoadQueue.scala 141:18:@4140.4]
  wire  entriesToCheck_1_7; // @[LoadQueue.scala 141:26:@4141.4]
  wire  _T_4706; // @[LoadQueue.scala 141:18:@4150.4]
  wire  entriesToCheck_2_0; // @[LoadQueue.scala 141:26:@4151.4]
  wire  _T_4708; // @[LoadQueue.scala 141:18:@4152.4]
  wire  entriesToCheck_2_1; // @[LoadQueue.scala 141:26:@4153.4]
  wire  _T_4710; // @[LoadQueue.scala 141:18:@4154.4]
  wire  entriesToCheck_2_2; // @[LoadQueue.scala 141:26:@4155.4]
  wire  _T_4712; // @[LoadQueue.scala 141:18:@4156.4]
  wire  entriesToCheck_2_3; // @[LoadQueue.scala 141:26:@4157.4]
  wire  _T_4714; // @[LoadQueue.scala 141:18:@4158.4]
  wire  entriesToCheck_2_4; // @[LoadQueue.scala 141:26:@4159.4]
  wire  _T_4716; // @[LoadQueue.scala 141:18:@4160.4]
  wire  entriesToCheck_2_5; // @[LoadQueue.scala 141:26:@4161.4]
  wire  _T_4718; // @[LoadQueue.scala 141:18:@4162.4]
  wire  entriesToCheck_2_6; // @[LoadQueue.scala 141:26:@4163.4]
  wire  _T_4720; // @[LoadQueue.scala 141:18:@4164.4]
  wire  entriesToCheck_2_7; // @[LoadQueue.scala 141:26:@4165.4]
  wire  _T_4722; // @[LoadQueue.scala 141:18:@4174.4]
  wire  entriesToCheck_3_0; // @[LoadQueue.scala 141:26:@4175.4]
  wire  _T_4724; // @[LoadQueue.scala 141:18:@4176.4]
  wire  entriesToCheck_3_1; // @[LoadQueue.scala 141:26:@4177.4]
  wire  _T_4726; // @[LoadQueue.scala 141:18:@4178.4]
  wire  entriesToCheck_3_2; // @[LoadQueue.scala 141:26:@4179.4]
  wire  _T_4728; // @[LoadQueue.scala 141:18:@4180.4]
  wire  entriesToCheck_3_3; // @[LoadQueue.scala 141:26:@4181.4]
  wire  _T_4730; // @[LoadQueue.scala 141:18:@4182.4]
  wire  entriesToCheck_3_4; // @[LoadQueue.scala 141:26:@4183.4]
  wire  _T_4732; // @[LoadQueue.scala 141:18:@4184.4]
  wire  entriesToCheck_3_5; // @[LoadQueue.scala 141:26:@4185.4]
  wire  _T_4734; // @[LoadQueue.scala 141:18:@4186.4]
  wire  entriesToCheck_3_6; // @[LoadQueue.scala 141:26:@4187.4]
  wire  _T_4736; // @[LoadQueue.scala 141:18:@4188.4]
  wire  entriesToCheck_3_7; // @[LoadQueue.scala 141:26:@4189.4]
  wire  _T_4738; // @[LoadQueue.scala 141:18:@4198.4]
  wire  entriesToCheck_4_0; // @[LoadQueue.scala 141:26:@4199.4]
  wire  _T_4740; // @[LoadQueue.scala 141:18:@4200.4]
  wire  entriesToCheck_4_1; // @[LoadQueue.scala 141:26:@4201.4]
  wire  _T_4742; // @[LoadQueue.scala 141:18:@4202.4]
  wire  entriesToCheck_4_2; // @[LoadQueue.scala 141:26:@4203.4]
  wire  _T_4744; // @[LoadQueue.scala 141:18:@4204.4]
  wire  entriesToCheck_4_3; // @[LoadQueue.scala 141:26:@4205.4]
  wire  _T_4746; // @[LoadQueue.scala 141:18:@4206.4]
  wire  entriesToCheck_4_4; // @[LoadQueue.scala 141:26:@4207.4]
  wire  _T_4748; // @[LoadQueue.scala 141:18:@4208.4]
  wire  entriesToCheck_4_5; // @[LoadQueue.scala 141:26:@4209.4]
  wire  _T_4750; // @[LoadQueue.scala 141:18:@4210.4]
  wire  entriesToCheck_4_6; // @[LoadQueue.scala 141:26:@4211.4]
  wire  _T_4752; // @[LoadQueue.scala 141:18:@4212.4]
  wire  entriesToCheck_4_7; // @[LoadQueue.scala 141:26:@4213.4]
  wire  _T_4754; // @[LoadQueue.scala 141:18:@4222.4]
  wire  entriesToCheck_5_0; // @[LoadQueue.scala 141:26:@4223.4]
  wire  _T_4756; // @[LoadQueue.scala 141:18:@4224.4]
  wire  entriesToCheck_5_1; // @[LoadQueue.scala 141:26:@4225.4]
  wire  _T_4758; // @[LoadQueue.scala 141:18:@4226.4]
  wire  entriesToCheck_5_2; // @[LoadQueue.scala 141:26:@4227.4]
  wire  _T_4760; // @[LoadQueue.scala 141:18:@4228.4]
  wire  entriesToCheck_5_3; // @[LoadQueue.scala 141:26:@4229.4]
  wire  _T_4762; // @[LoadQueue.scala 141:18:@4230.4]
  wire  entriesToCheck_5_4; // @[LoadQueue.scala 141:26:@4231.4]
  wire  _T_4764; // @[LoadQueue.scala 141:18:@4232.4]
  wire  entriesToCheck_5_5; // @[LoadQueue.scala 141:26:@4233.4]
  wire  _T_4766; // @[LoadQueue.scala 141:18:@4234.4]
  wire  entriesToCheck_5_6; // @[LoadQueue.scala 141:26:@4235.4]
  wire  _T_4768; // @[LoadQueue.scala 141:18:@4236.4]
  wire  entriesToCheck_5_7; // @[LoadQueue.scala 141:26:@4237.4]
  wire  _T_4770; // @[LoadQueue.scala 141:18:@4246.4]
  wire  entriesToCheck_6_0; // @[LoadQueue.scala 141:26:@4247.4]
  wire  _T_4772; // @[LoadQueue.scala 141:18:@4248.4]
  wire  entriesToCheck_6_1; // @[LoadQueue.scala 141:26:@4249.4]
  wire  _T_4774; // @[LoadQueue.scala 141:18:@4250.4]
  wire  entriesToCheck_6_2; // @[LoadQueue.scala 141:26:@4251.4]
  wire  _T_4776; // @[LoadQueue.scala 141:18:@4252.4]
  wire  entriesToCheck_6_3; // @[LoadQueue.scala 141:26:@4253.4]
  wire  _T_4778; // @[LoadQueue.scala 141:18:@4254.4]
  wire  entriesToCheck_6_4; // @[LoadQueue.scala 141:26:@4255.4]
  wire  _T_4780; // @[LoadQueue.scala 141:18:@4256.4]
  wire  entriesToCheck_6_5; // @[LoadQueue.scala 141:26:@4257.4]
  wire  _T_4782; // @[LoadQueue.scala 141:18:@4258.4]
  wire  entriesToCheck_6_6; // @[LoadQueue.scala 141:26:@4259.4]
  wire  _T_4784; // @[LoadQueue.scala 141:18:@4260.4]
  wire  entriesToCheck_6_7; // @[LoadQueue.scala 141:26:@4261.4]
  wire  _T_4786; // @[LoadQueue.scala 141:18:@4270.4]
  wire  entriesToCheck_7_0; // @[LoadQueue.scala 141:26:@4271.4]
  wire  _T_4788; // @[LoadQueue.scala 141:18:@4272.4]
  wire  entriesToCheck_7_1; // @[LoadQueue.scala 141:26:@4273.4]
  wire  _T_4790; // @[LoadQueue.scala 141:18:@4274.4]
  wire  entriesToCheck_7_2; // @[LoadQueue.scala 141:26:@4275.4]
  wire  _T_4792; // @[LoadQueue.scala 141:18:@4276.4]
  wire  entriesToCheck_7_3; // @[LoadQueue.scala 141:26:@4277.4]
  wire  _T_4794; // @[LoadQueue.scala 141:18:@4278.4]
  wire  entriesToCheck_7_4; // @[LoadQueue.scala 141:26:@4279.4]
  wire  _T_4796; // @[LoadQueue.scala 141:18:@4280.4]
  wire  entriesToCheck_7_5; // @[LoadQueue.scala 141:26:@4281.4]
  wire  _T_4798; // @[LoadQueue.scala 141:18:@4282.4]
  wire  entriesToCheck_7_6; // @[LoadQueue.scala 141:26:@4283.4]
  wire  _T_4800; // @[LoadQueue.scala 141:18:@4284.4]
  wire  entriesToCheck_7_7; // @[LoadQueue.scala 141:26:@4285.4]
  wire  _T_5168; // @[LoadQueue.scala 151:92:@4295.4]
  wire  _T_5169; // @[LoadQueue.scala 152:41:@4296.4]
  wire  _T_5170; // @[LoadQueue.scala 153:30:@4297.4]
  wire  conflict_0_0; // @[LoadQueue.scala 152:68:@4298.4]
  wire  _T_5172; // @[LoadQueue.scala 151:92:@4300.4]
  wire  _T_5173; // @[LoadQueue.scala 152:41:@4301.4]
  wire  _T_5174; // @[LoadQueue.scala 153:30:@4302.4]
  wire  conflict_0_1; // @[LoadQueue.scala 152:68:@4303.4]
  wire  _T_5176; // @[LoadQueue.scala 151:92:@4305.4]
  wire  _T_5177; // @[LoadQueue.scala 152:41:@4306.4]
  wire  _T_5178; // @[LoadQueue.scala 153:30:@4307.4]
  wire  conflict_0_2; // @[LoadQueue.scala 152:68:@4308.4]
  wire  _T_5180; // @[LoadQueue.scala 151:92:@4310.4]
  wire  _T_5181; // @[LoadQueue.scala 152:41:@4311.4]
  wire  _T_5182; // @[LoadQueue.scala 153:30:@4312.4]
  wire  conflict_0_3; // @[LoadQueue.scala 152:68:@4313.4]
  wire  _T_5184; // @[LoadQueue.scala 151:92:@4315.4]
  wire  _T_5185; // @[LoadQueue.scala 152:41:@4316.4]
  wire  _T_5186; // @[LoadQueue.scala 153:30:@4317.4]
  wire  conflict_0_4; // @[LoadQueue.scala 152:68:@4318.4]
  wire  _T_5188; // @[LoadQueue.scala 151:92:@4320.4]
  wire  _T_5189; // @[LoadQueue.scala 152:41:@4321.4]
  wire  _T_5190; // @[LoadQueue.scala 153:30:@4322.4]
  wire  conflict_0_5; // @[LoadQueue.scala 152:68:@4323.4]
  wire  _T_5192; // @[LoadQueue.scala 151:92:@4325.4]
  wire  _T_5193; // @[LoadQueue.scala 152:41:@4326.4]
  wire  _T_5194; // @[LoadQueue.scala 153:30:@4327.4]
  wire  conflict_0_6; // @[LoadQueue.scala 152:68:@4328.4]
  wire  _T_5196; // @[LoadQueue.scala 151:92:@4330.4]
  wire  _T_5197; // @[LoadQueue.scala 152:41:@4331.4]
  wire  _T_5198; // @[LoadQueue.scala 153:30:@4332.4]
  wire  conflict_0_7; // @[LoadQueue.scala 152:68:@4333.4]
  wire  _T_5200; // @[LoadQueue.scala 151:92:@4335.4]
  wire  _T_5201; // @[LoadQueue.scala 152:41:@4336.4]
  wire  _T_5202; // @[LoadQueue.scala 153:30:@4337.4]
  wire  conflict_1_0; // @[LoadQueue.scala 152:68:@4338.4]
  wire  _T_5204; // @[LoadQueue.scala 151:92:@4340.4]
  wire  _T_5205; // @[LoadQueue.scala 152:41:@4341.4]
  wire  _T_5206; // @[LoadQueue.scala 153:30:@4342.4]
  wire  conflict_1_1; // @[LoadQueue.scala 152:68:@4343.4]
  wire  _T_5208; // @[LoadQueue.scala 151:92:@4345.4]
  wire  _T_5209; // @[LoadQueue.scala 152:41:@4346.4]
  wire  _T_5210; // @[LoadQueue.scala 153:30:@4347.4]
  wire  conflict_1_2; // @[LoadQueue.scala 152:68:@4348.4]
  wire  _T_5212; // @[LoadQueue.scala 151:92:@4350.4]
  wire  _T_5213; // @[LoadQueue.scala 152:41:@4351.4]
  wire  _T_5214; // @[LoadQueue.scala 153:30:@4352.4]
  wire  conflict_1_3; // @[LoadQueue.scala 152:68:@4353.4]
  wire  _T_5216; // @[LoadQueue.scala 151:92:@4355.4]
  wire  _T_5217; // @[LoadQueue.scala 152:41:@4356.4]
  wire  _T_5218; // @[LoadQueue.scala 153:30:@4357.4]
  wire  conflict_1_4; // @[LoadQueue.scala 152:68:@4358.4]
  wire  _T_5220; // @[LoadQueue.scala 151:92:@4360.4]
  wire  _T_5221; // @[LoadQueue.scala 152:41:@4361.4]
  wire  _T_5222; // @[LoadQueue.scala 153:30:@4362.4]
  wire  conflict_1_5; // @[LoadQueue.scala 152:68:@4363.4]
  wire  _T_5224; // @[LoadQueue.scala 151:92:@4365.4]
  wire  _T_5225; // @[LoadQueue.scala 152:41:@4366.4]
  wire  _T_5226; // @[LoadQueue.scala 153:30:@4367.4]
  wire  conflict_1_6; // @[LoadQueue.scala 152:68:@4368.4]
  wire  _T_5228; // @[LoadQueue.scala 151:92:@4370.4]
  wire  _T_5229; // @[LoadQueue.scala 152:41:@4371.4]
  wire  _T_5230; // @[LoadQueue.scala 153:30:@4372.4]
  wire  conflict_1_7; // @[LoadQueue.scala 152:68:@4373.4]
  wire  _T_5232; // @[LoadQueue.scala 151:92:@4375.4]
  wire  _T_5233; // @[LoadQueue.scala 152:41:@4376.4]
  wire  _T_5234; // @[LoadQueue.scala 153:30:@4377.4]
  wire  conflict_2_0; // @[LoadQueue.scala 152:68:@4378.4]
  wire  _T_5236; // @[LoadQueue.scala 151:92:@4380.4]
  wire  _T_5237; // @[LoadQueue.scala 152:41:@4381.4]
  wire  _T_5238; // @[LoadQueue.scala 153:30:@4382.4]
  wire  conflict_2_1; // @[LoadQueue.scala 152:68:@4383.4]
  wire  _T_5240; // @[LoadQueue.scala 151:92:@4385.4]
  wire  _T_5241; // @[LoadQueue.scala 152:41:@4386.4]
  wire  _T_5242; // @[LoadQueue.scala 153:30:@4387.4]
  wire  conflict_2_2; // @[LoadQueue.scala 152:68:@4388.4]
  wire  _T_5244; // @[LoadQueue.scala 151:92:@4390.4]
  wire  _T_5245; // @[LoadQueue.scala 152:41:@4391.4]
  wire  _T_5246; // @[LoadQueue.scala 153:30:@4392.4]
  wire  conflict_2_3; // @[LoadQueue.scala 152:68:@4393.4]
  wire  _T_5248; // @[LoadQueue.scala 151:92:@4395.4]
  wire  _T_5249; // @[LoadQueue.scala 152:41:@4396.4]
  wire  _T_5250; // @[LoadQueue.scala 153:30:@4397.4]
  wire  conflict_2_4; // @[LoadQueue.scala 152:68:@4398.4]
  wire  _T_5252; // @[LoadQueue.scala 151:92:@4400.4]
  wire  _T_5253; // @[LoadQueue.scala 152:41:@4401.4]
  wire  _T_5254; // @[LoadQueue.scala 153:30:@4402.4]
  wire  conflict_2_5; // @[LoadQueue.scala 152:68:@4403.4]
  wire  _T_5256; // @[LoadQueue.scala 151:92:@4405.4]
  wire  _T_5257; // @[LoadQueue.scala 152:41:@4406.4]
  wire  _T_5258; // @[LoadQueue.scala 153:30:@4407.4]
  wire  conflict_2_6; // @[LoadQueue.scala 152:68:@4408.4]
  wire  _T_5260; // @[LoadQueue.scala 151:92:@4410.4]
  wire  _T_5261; // @[LoadQueue.scala 152:41:@4411.4]
  wire  _T_5262; // @[LoadQueue.scala 153:30:@4412.4]
  wire  conflict_2_7; // @[LoadQueue.scala 152:68:@4413.4]
  wire  _T_5264; // @[LoadQueue.scala 151:92:@4415.4]
  wire  _T_5265; // @[LoadQueue.scala 152:41:@4416.4]
  wire  _T_5266; // @[LoadQueue.scala 153:30:@4417.4]
  wire  conflict_3_0; // @[LoadQueue.scala 152:68:@4418.4]
  wire  _T_5268; // @[LoadQueue.scala 151:92:@4420.4]
  wire  _T_5269; // @[LoadQueue.scala 152:41:@4421.4]
  wire  _T_5270; // @[LoadQueue.scala 153:30:@4422.4]
  wire  conflict_3_1; // @[LoadQueue.scala 152:68:@4423.4]
  wire  _T_5272; // @[LoadQueue.scala 151:92:@4425.4]
  wire  _T_5273; // @[LoadQueue.scala 152:41:@4426.4]
  wire  _T_5274; // @[LoadQueue.scala 153:30:@4427.4]
  wire  conflict_3_2; // @[LoadQueue.scala 152:68:@4428.4]
  wire  _T_5276; // @[LoadQueue.scala 151:92:@4430.4]
  wire  _T_5277; // @[LoadQueue.scala 152:41:@4431.4]
  wire  _T_5278; // @[LoadQueue.scala 153:30:@4432.4]
  wire  conflict_3_3; // @[LoadQueue.scala 152:68:@4433.4]
  wire  _T_5280; // @[LoadQueue.scala 151:92:@4435.4]
  wire  _T_5281; // @[LoadQueue.scala 152:41:@4436.4]
  wire  _T_5282; // @[LoadQueue.scala 153:30:@4437.4]
  wire  conflict_3_4; // @[LoadQueue.scala 152:68:@4438.4]
  wire  _T_5284; // @[LoadQueue.scala 151:92:@4440.4]
  wire  _T_5285; // @[LoadQueue.scala 152:41:@4441.4]
  wire  _T_5286; // @[LoadQueue.scala 153:30:@4442.4]
  wire  conflict_3_5; // @[LoadQueue.scala 152:68:@4443.4]
  wire  _T_5288; // @[LoadQueue.scala 151:92:@4445.4]
  wire  _T_5289; // @[LoadQueue.scala 152:41:@4446.4]
  wire  _T_5290; // @[LoadQueue.scala 153:30:@4447.4]
  wire  conflict_3_6; // @[LoadQueue.scala 152:68:@4448.4]
  wire  _T_5292; // @[LoadQueue.scala 151:92:@4450.4]
  wire  _T_5293; // @[LoadQueue.scala 152:41:@4451.4]
  wire  _T_5294; // @[LoadQueue.scala 153:30:@4452.4]
  wire  conflict_3_7; // @[LoadQueue.scala 152:68:@4453.4]
  wire  _T_5296; // @[LoadQueue.scala 151:92:@4455.4]
  wire  _T_5297; // @[LoadQueue.scala 152:41:@4456.4]
  wire  _T_5298; // @[LoadQueue.scala 153:30:@4457.4]
  wire  conflict_4_0; // @[LoadQueue.scala 152:68:@4458.4]
  wire  _T_5300; // @[LoadQueue.scala 151:92:@4460.4]
  wire  _T_5301; // @[LoadQueue.scala 152:41:@4461.4]
  wire  _T_5302; // @[LoadQueue.scala 153:30:@4462.4]
  wire  conflict_4_1; // @[LoadQueue.scala 152:68:@4463.4]
  wire  _T_5304; // @[LoadQueue.scala 151:92:@4465.4]
  wire  _T_5305; // @[LoadQueue.scala 152:41:@4466.4]
  wire  _T_5306; // @[LoadQueue.scala 153:30:@4467.4]
  wire  conflict_4_2; // @[LoadQueue.scala 152:68:@4468.4]
  wire  _T_5308; // @[LoadQueue.scala 151:92:@4470.4]
  wire  _T_5309; // @[LoadQueue.scala 152:41:@4471.4]
  wire  _T_5310; // @[LoadQueue.scala 153:30:@4472.4]
  wire  conflict_4_3; // @[LoadQueue.scala 152:68:@4473.4]
  wire  _T_5312; // @[LoadQueue.scala 151:92:@4475.4]
  wire  _T_5313; // @[LoadQueue.scala 152:41:@4476.4]
  wire  _T_5314; // @[LoadQueue.scala 153:30:@4477.4]
  wire  conflict_4_4; // @[LoadQueue.scala 152:68:@4478.4]
  wire  _T_5316; // @[LoadQueue.scala 151:92:@4480.4]
  wire  _T_5317; // @[LoadQueue.scala 152:41:@4481.4]
  wire  _T_5318; // @[LoadQueue.scala 153:30:@4482.4]
  wire  conflict_4_5; // @[LoadQueue.scala 152:68:@4483.4]
  wire  _T_5320; // @[LoadQueue.scala 151:92:@4485.4]
  wire  _T_5321; // @[LoadQueue.scala 152:41:@4486.4]
  wire  _T_5322; // @[LoadQueue.scala 153:30:@4487.4]
  wire  conflict_4_6; // @[LoadQueue.scala 152:68:@4488.4]
  wire  _T_5324; // @[LoadQueue.scala 151:92:@4490.4]
  wire  _T_5325; // @[LoadQueue.scala 152:41:@4491.4]
  wire  _T_5326; // @[LoadQueue.scala 153:30:@4492.4]
  wire  conflict_4_7; // @[LoadQueue.scala 152:68:@4493.4]
  wire  _T_5328; // @[LoadQueue.scala 151:92:@4495.4]
  wire  _T_5329; // @[LoadQueue.scala 152:41:@4496.4]
  wire  _T_5330; // @[LoadQueue.scala 153:30:@4497.4]
  wire  conflict_5_0; // @[LoadQueue.scala 152:68:@4498.4]
  wire  _T_5332; // @[LoadQueue.scala 151:92:@4500.4]
  wire  _T_5333; // @[LoadQueue.scala 152:41:@4501.4]
  wire  _T_5334; // @[LoadQueue.scala 153:30:@4502.4]
  wire  conflict_5_1; // @[LoadQueue.scala 152:68:@4503.4]
  wire  _T_5336; // @[LoadQueue.scala 151:92:@4505.4]
  wire  _T_5337; // @[LoadQueue.scala 152:41:@4506.4]
  wire  _T_5338; // @[LoadQueue.scala 153:30:@4507.4]
  wire  conflict_5_2; // @[LoadQueue.scala 152:68:@4508.4]
  wire  _T_5340; // @[LoadQueue.scala 151:92:@4510.4]
  wire  _T_5341; // @[LoadQueue.scala 152:41:@4511.4]
  wire  _T_5342; // @[LoadQueue.scala 153:30:@4512.4]
  wire  conflict_5_3; // @[LoadQueue.scala 152:68:@4513.4]
  wire  _T_5344; // @[LoadQueue.scala 151:92:@4515.4]
  wire  _T_5345; // @[LoadQueue.scala 152:41:@4516.4]
  wire  _T_5346; // @[LoadQueue.scala 153:30:@4517.4]
  wire  conflict_5_4; // @[LoadQueue.scala 152:68:@4518.4]
  wire  _T_5348; // @[LoadQueue.scala 151:92:@4520.4]
  wire  _T_5349; // @[LoadQueue.scala 152:41:@4521.4]
  wire  _T_5350; // @[LoadQueue.scala 153:30:@4522.4]
  wire  conflict_5_5; // @[LoadQueue.scala 152:68:@4523.4]
  wire  _T_5352; // @[LoadQueue.scala 151:92:@4525.4]
  wire  _T_5353; // @[LoadQueue.scala 152:41:@4526.4]
  wire  _T_5354; // @[LoadQueue.scala 153:30:@4527.4]
  wire  conflict_5_6; // @[LoadQueue.scala 152:68:@4528.4]
  wire  _T_5356; // @[LoadQueue.scala 151:92:@4530.4]
  wire  _T_5357; // @[LoadQueue.scala 152:41:@4531.4]
  wire  _T_5358; // @[LoadQueue.scala 153:30:@4532.4]
  wire  conflict_5_7; // @[LoadQueue.scala 152:68:@4533.4]
  wire  _T_5360; // @[LoadQueue.scala 151:92:@4535.4]
  wire  _T_5361; // @[LoadQueue.scala 152:41:@4536.4]
  wire  _T_5362; // @[LoadQueue.scala 153:30:@4537.4]
  wire  conflict_6_0; // @[LoadQueue.scala 152:68:@4538.4]
  wire  _T_5364; // @[LoadQueue.scala 151:92:@4540.4]
  wire  _T_5365; // @[LoadQueue.scala 152:41:@4541.4]
  wire  _T_5366; // @[LoadQueue.scala 153:30:@4542.4]
  wire  conflict_6_1; // @[LoadQueue.scala 152:68:@4543.4]
  wire  _T_5368; // @[LoadQueue.scala 151:92:@4545.4]
  wire  _T_5369; // @[LoadQueue.scala 152:41:@4546.4]
  wire  _T_5370; // @[LoadQueue.scala 153:30:@4547.4]
  wire  conflict_6_2; // @[LoadQueue.scala 152:68:@4548.4]
  wire  _T_5372; // @[LoadQueue.scala 151:92:@4550.4]
  wire  _T_5373; // @[LoadQueue.scala 152:41:@4551.4]
  wire  _T_5374; // @[LoadQueue.scala 153:30:@4552.4]
  wire  conflict_6_3; // @[LoadQueue.scala 152:68:@4553.4]
  wire  _T_5376; // @[LoadQueue.scala 151:92:@4555.4]
  wire  _T_5377; // @[LoadQueue.scala 152:41:@4556.4]
  wire  _T_5378; // @[LoadQueue.scala 153:30:@4557.4]
  wire  conflict_6_4; // @[LoadQueue.scala 152:68:@4558.4]
  wire  _T_5380; // @[LoadQueue.scala 151:92:@4560.4]
  wire  _T_5381; // @[LoadQueue.scala 152:41:@4561.4]
  wire  _T_5382; // @[LoadQueue.scala 153:30:@4562.4]
  wire  conflict_6_5; // @[LoadQueue.scala 152:68:@4563.4]
  wire  _T_5384; // @[LoadQueue.scala 151:92:@4565.4]
  wire  _T_5385; // @[LoadQueue.scala 152:41:@4566.4]
  wire  _T_5386; // @[LoadQueue.scala 153:30:@4567.4]
  wire  conflict_6_6; // @[LoadQueue.scala 152:68:@4568.4]
  wire  _T_5388; // @[LoadQueue.scala 151:92:@4570.4]
  wire  _T_5389; // @[LoadQueue.scala 152:41:@4571.4]
  wire  _T_5390; // @[LoadQueue.scala 153:30:@4572.4]
  wire  conflict_6_7; // @[LoadQueue.scala 152:68:@4573.4]
  wire  _T_5392; // @[LoadQueue.scala 151:92:@4575.4]
  wire  _T_5393; // @[LoadQueue.scala 152:41:@4576.4]
  wire  _T_5394; // @[LoadQueue.scala 153:30:@4577.4]
  wire  conflict_7_0; // @[LoadQueue.scala 152:68:@4578.4]
  wire  _T_5396; // @[LoadQueue.scala 151:92:@4580.4]
  wire  _T_5397; // @[LoadQueue.scala 152:41:@4581.4]
  wire  _T_5398; // @[LoadQueue.scala 153:30:@4582.4]
  wire  conflict_7_1; // @[LoadQueue.scala 152:68:@4583.4]
  wire  _T_5400; // @[LoadQueue.scala 151:92:@4585.4]
  wire  _T_5401; // @[LoadQueue.scala 152:41:@4586.4]
  wire  _T_5402; // @[LoadQueue.scala 153:30:@4587.4]
  wire  conflict_7_2; // @[LoadQueue.scala 152:68:@4588.4]
  wire  _T_5404; // @[LoadQueue.scala 151:92:@4590.4]
  wire  _T_5405; // @[LoadQueue.scala 152:41:@4591.4]
  wire  _T_5406; // @[LoadQueue.scala 153:30:@4592.4]
  wire  conflict_7_3; // @[LoadQueue.scala 152:68:@4593.4]
  wire  _T_5408; // @[LoadQueue.scala 151:92:@4595.4]
  wire  _T_5409; // @[LoadQueue.scala 152:41:@4596.4]
  wire  _T_5410; // @[LoadQueue.scala 153:30:@4597.4]
  wire  conflict_7_4; // @[LoadQueue.scala 152:68:@4598.4]
  wire  _T_5412; // @[LoadQueue.scala 151:92:@4600.4]
  wire  _T_5413; // @[LoadQueue.scala 152:41:@4601.4]
  wire  _T_5414; // @[LoadQueue.scala 153:30:@4602.4]
  wire  conflict_7_5; // @[LoadQueue.scala 152:68:@4603.4]
  wire  _T_5416; // @[LoadQueue.scala 151:92:@4605.4]
  wire  _T_5417; // @[LoadQueue.scala 152:41:@4606.4]
  wire  _T_5418; // @[LoadQueue.scala 153:30:@4607.4]
  wire  conflict_7_6; // @[LoadQueue.scala 152:68:@4608.4]
  wire  _T_5420; // @[LoadQueue.scala 151:92:@4610.4]
  wire  _T_5421; // @[LoadQueue.scala 152:41:@4611.4]
  wire  _T_5422; // @[LoadQueue.scala 153:30:@4612.4]
  wire  conflict_7_7; // @[LoadQueue.scala 152:68:@4613.4]
  wire  _T_5791; // @[LoadQueue.scala 163:13:@4616.4]
  wire  storeAddrNotKnownFlags_0_0; // @[LoadQueue.scala 163:19:@4617.4]
  wire  _T_5794; // @[LoadQueue.scala 163:13:@4618.4]
  wire  storeAddrNotKnownFlags_0_1; // @[LoadQueue.scala 163:19:@4619.4]
  wire  _T_5797; // @[LoadQueue.scala 163:13:@4620.4]
  wire  storeAddrNotKnownFlags_0_2; // @[LoadQueue.scala 163:19:@4621.4]
  wire  _T_5800; // @[LoadQueue.scala 163:13:@4622.4]
  wire  storeAddrNotKnownFlags_0_3; // @[LoadQueue.scala 163:19:@4623.4]
  wire  _T_5803; // @[LoadQueue.scala 163:13:@4624.4]
  wire  storeAddrNotKnownFlags_0_4; // @[LoadQueue.scala 163:19:@4625.4]
  wire  _T_5806; // @[LoadQueue.scala 163:13:@4626.4]
  wire  storeAddrNotKnownFlags_0_5; // @[LoadQueue.scala 163:19:@4627.4]
  wire  _T_5809; // @[LoadQueue.scala 163:13:@4628.4]
  wire  storeAddrNotKnownFlags_0_6; // @[LoadQueue.scala 163:19:@4629.4]
  wire  _T_5812; // @[LoadQueue.scala 163:13:@4630.4]
  wire  storeAddrNotKnownFlags_0_7; // @[LoadQueue.scala 163:19:@4631.4]
  wire  storeAddrNotKnownFlags_1_0; // @[LoadQueue.scala 163:19:@4641.4]
  wire  storeAddrNotKnownFlags_1_1; // @[LoadQueue.scala 163:19:@4643.4]
  wire  storeAddrNotKnownFlags_1_2; // @[LoadQueue.scala 163:19:@4645.4]
  wire  storeAddrNotKnownFlags_1_3; // @[LoadQueue.scala 163:19:@4647.4]
  wire  storeAddrNotKnownFlags_1_4; // @[LoadQueue.scala 163:19:@4649.4]
  wire  storeAddrNotKnownFlags_1_5; // @[LoadQueue.scala 163:19:@4651.4]
  wire  storeAddrNotKnownFlags_1_6; // @[LoadQueue.scala 163:19:@4653.4]
  wire  storeAddrNotKnownFlags_1_7; // @[LoadQueue.scala 163:19:@4655.4]
  wire  storeAddrNotKnownFlags_2_0; // @[LoadQueue.scala 163:19:@4665.4]
  wire  storeAddrNotKnownFlags_2_1; // @[LoadQueue.scala 163:19:@4667.4]
  wire  storeAddrNotKnownFlags_2_2; // @[LoadQueue.scala 163:19:@4669.4]
  wire  storeAddrNotKnownFlags_2_3; // @[LoadQueue.scala 163:19:@4671.4]
  wire  storeAddrNotKnownFlags_2_4; // @[LoadQueue.scala 163:19:@4673.4]
  wire  storeAddrNotKnownFlags_2_5; // @[LoadQueue.scala 163:19:@4675.4]
  wire  storeAddrNotKnownFlags_2_6; // @[LoadQueue.scala 163:19:@4677.4]
  wire  storeAddrNotKnownFlags_2_7; // @[LoadQueue.scala 163:19:@4679.4]
  wire  storeAddrNotKnownFlags_3_0; // @[LoadQueue.scala 163:19:@4689.4]
  wire  storeAddrNotKnownFlags_3_1; // @[LoadQueue.scala 163:19:@4691.4]
  wire  storeAddrNotKnownFlags_3_2; // @[LoadQueue.scala 163:19:@4693.4]
  wire  storeAddrNotKnownFlags_3_3; // @[LoadQueue.scala 163:19:@4695.4]
  wire  storeAddrNotKnownFlags_3_4; // @[LoadQueue.scala 163:19:@4697.4]
  wire  storeAddrNotKnownFlags_3_5; // @[LoadQueue.scala 163:19:@4699.4]
  wire  storeAddrNotKnownFlags_3_6; // @[LoadQueue.scala 163:19:@4701.4]
  wire  storeAddrNotKnownFlags_3_7; // @[LoadQueue.scala 163:19:@4703.4]
  wire  storeAddrNotKnownFlags_4_0; // @[LoadQueue.scala 163:19:@4713.4]
  wire  storeAddrNotKnownFlags_4_1; // @[LoadQueue.scala 163:19:@4715.4]
  wire  storeAddrNotKnownFlags_4_2; // @[LoadQueue.scala 163:19:@4717.4]
  wire  storeAddrNotKnownFlags_4_3; // @[LoadQueue.scala 163:19:@4719.4]
  wire  storeAddrNotKnownFlags_4_4; // @[LoadQueue.scala 163:19:@4721.4]
  wire  storeAddrNotKnownFlags_4_5; // @[LoadQueue.scala 163:19:@4723.4]
  wire  storeAddrNotKnownFlags_4_6; // @[LoadQueue.scala 163:19:@4725.4]
  wire  storeAddrNotKnownFlags_4_7; // @[LoadQueue.scala 163:19:@4727.4]
  wire  storeAddrNotKnownFlags_5_0; // @[LoadQueue.scala 163:19:@4737.4]
  wire  storeAddrNotKnownFlags_5_1; // @[LoadQueue.scala 163:19:@4739.4]
  wire  storeAddrNotKnownFlags_5_2; // @[LoadQueue.scala 163:19:@4741.4]
  wire  storeAddrNotKnownFlags_5_3; // @[LoadQueue.scala 163:19:@4743.4]
  wire  storeAddrNotKnownFlags_5_4; // @[LoadQueue.scala 163:19:@4745.4]
  wire  storeAddrNotKnownFlags_5_5; // @[LoadQueue.scala 163:19:@4747.4]
  wire  storeAddrNotKnownFlags_5_6; // @[LoadQueue.scala 163:19:@4749.4]
  wire  storeAddrNotKnownFlags_5_7; // @[LoadQueue.scala 163:19:@4751.4]
  wire  storeAddrNotKnownFlags_6_0; // @[LoadQueue.scala 163:19:@4761.4]
  wire  storeAddrNotKnownFlags_6_1; // @[LoadQueue.scala 163:19:@4763.4]
  wire  storeAddrNotKnownFlags_6_2; // @[LoadQueue.scala 163:19:@4765.4]
  wire  storeAddrNotKnownFlags_6_3; // @[LoadQueue.scala 163:19:@4767.4]
  wire  storeAddrNotKnownFlags_6_4; // @[LoadQueue.scala 163:19:@4769.4]
  wire  storeAddrNotKnownFlags_6_5; // @[LoadQueue.scala 163:19:@4771.4]
  wire  storeAddrNotKnownFlags_6_6; // @[LoadQueue.scala 163:19:@4773.4]
  wire  storeAddrNotKnownFlags_6_7; // @[LoadQueue.scala 163:19:@4775.4]
  wire  storeAddrNotKnownFlags_7_0; // @[LoadQueue.scala 163:19:@4785.4]
  wire  storeAddrNotKnownFlags_7_1; // @[LoadQueue.scala 163:19:@4787.4]
  wire  storeAddrNotKnownFlags_7_2; // @[LoadQueue.scala 163:19:@4789.4]
  wire  storeAddrNotKnownFlags_7_3; // @[LoadQueue.scala 163:19:@4791.4]
  wire  storeAddrNotKnownFlags_7_4; // @[LoadQueue.scala 163:19:@4793.4]
  wire  storeAddrNotKnownFlags_7_5; // @[LoadQueue.scala 163:19:@4795.4]
  wire  storeAddrNotKnownFlags_7_6; // @[LoadQueue.scala 163:19:@4797.4]
  wire  storeAddrNotKnownFlags_7_7; // @[LoadQueue.scala 163:19:@4799.4]
  wire [7:0] _T_6146; // @[Mux.scala 19:72:@4906.4]
  wire [7:0] _T_6148; // @[Mux.scala 19:72:@4907.4]
  wire [7:0] _T_6155; // @[Mux.scala 19:72:@4914.4]
  wire [7:0] _T_6157; // @[Mux.scala 19:72:@4915.4]
  wire [7:0] _T_6164; // @[Mux.scala 19:72:@4922.4]
  wire [7:0] _T_6166; // @[Mux.scala 19:72:@4923.4]
  wire [7:0] _T_6173; // @[Mux.scala 19:72:@4930.4]
  wire [7:0] _T_6175; // @[Mux.scala 19:72:@4931.4]
  wire [7:0] _T_6182; // @[Mux.scala 19:72:@4938.4]
  wire [7:0] _T_6184; // @[Mux.scala 19:72:@4939.4]
  wire [7:0] _T_6191; // @[Mux.scala 19:72:@4946.4]
  wire [7:0] _T_6193; // @[Mux.scala 19:72:@4947.4]
  wire [7:0] _T_6200; // @[Mux.scala 19:72:@4954.4]
  wire [7:0] _T_6202; // @[Mux.scala 19:72:@4955.4]
  wire [7:0] _T_6209; // @[Mux.scala 19:72:@4962.4]
  wire [7:0] _T_6211; // @[Mux.scala 19:72:@4963.4]
  wire [7:0] _T_6212; // @[Mux.scala 19:72:@4964.4]
  wire [7:0] _T_6213; // @[Mux.scala 19:72:@4965.4]
  wire [7:0] _T_6214; // @[Mux.scala 19:72:@4966.4]
  wire [7:0] _T_6215; // @[Mux.scala 19:72:@4967.4]
  wire [7:0] _T_6216; // @[Mux.scala 19:72:@4968.4]
  wire [7:0] _T_6217; // @[Mux.scala 19:72:@4969.4]
  wire [7:0] _T_6218; // @[Mux.scala 19:72:@4970.4]
  wire [7:0] _T_6460; // @[Mux.scala 19:72:@5088.4]
  wire [7:0] _T_6462; // @[Mux.scala 19:72:@5089.4]
  wire [7:0] _T_6469; // @[Mux.scala 19:72:@5096.4]
  wire [7:0] _T_6471; // @[Mux.scala 19:72:@5097.4]
  wire [7:0] _T_6478; // @[Mux.scala 19:72:@5104.4]
  wire [7:0] _T_6480; // @[Mux.scala 19:72:@5105.4]
  wire [7:0] _T_6487; // @[Mux.scala 19:72:@5112.4]
  wire [7:0] _T_6489; // @[Mux.scala 19:72:@5113.4]
  wire [7:0] _T_6496; // @[Mux.scala 19:72:@5120.4]
  wire [7:0] _T_6498; // @[Mux.scala 19:72:@5121.4]
  wire [7:0] _T_6505; // @[Mux.scala 19:72:@5128.4]
  wire [7:0] _T_6507; // @[Mux.scala 19:72:@5129.4]
  wire [7:0] _T_6514; // @[Mux.scala 19:72:@5136.4]
  wire [7:0] _T_6516; // @[Mux.scala 19:72:@5137.4]
  wire [7:0] _T_6523; // @[Mux.scala 19:72:@5144.4]
  wire [7:0] _T_6525; // @[Mux.scala 19:72:@5145.4]
  wire [7:0] _T_6526; // @[Mux.scala 19:72:@5146.4]
  wire [7:0] _T_6527; // @[Mux.scala 19:72:@5147.4]
  wire [7:0] _T_6528; // @[Mux.scala 19:72:@5148.4]
  wire [7:0] _T_6529; // @[Mux.scala 19:72:@5149.4]
  wire [7:0] _T_6530; // @[Mux.scala 19:72:@5150.4]
  wire [7:0] _T_6531; // @[Mux.scala 19:72:@5151.4]
  wire [7:0] _T_6532; // @[Mux.scala 19:72:@5152.4]
  wire [7:0] _T_6774; // @[Mux.scala 19:72:@5270.4]
  wire [7:0] _T_6776; // @[Mux.scala 19:72:@5271.4]
  wire [7:0] _T_6783; // @[Mux.scala 19:72:@5278.4]
  wire [7:0] _T_6785; // @[Mux.scala 19:72:@5279.4]
  wire [7:0] _T_6792; // @[Mux.scala 19:72:@5286.4]
  wire [7:0] _T_6794; // @[Mux.scala 19:72:@5287.4]
  wire [7:0] _T_6801; // @[Mux.scala 19:72:@5294.4]
  wire [7:0] _T_6803; // @[Mux.scala 19:72:@5295.4]
  wire [7:0] _T_6810; // @[Mux.scala 19:72:@5302.4]
  wire [7:0] _T_6812; // @[Mux.scala 19:72:@5303.4]
  wire [7:0] _T_6819; // @[Mux.scala 19:72:@5310.4]
  wire [7:0] _T_6821; // @[Mux.scala 19:72:@5311.4]
  wire [7:0] _T_6828; // @[Mux.scala 19:72:@5318.4]
  wire [7:0] _T_6830; // @[Mux.scala 19:72:@5319.4]
  wire [7:0] _T_6837; // @[Mux.scala 19:72:@5326.4]
  wire [7:0] _T_6839; // @[Mux.scala 19:72:@5327.4]
  wire [7:0] _T_6840; // @[Mux.scala 19:72:@5328.4]
  wire [7:0] _T_6841; // @[Mux.scala 19:72:@5329.4]
  wire [7:0] _T_6842; // @[Mux.scala 19:72:@5330.4]
  wire [7:0] _T_6843; // @[Mux.scala 19:72:@5331.4]
  wire [7:0] _T_6844; // @[Mux.scala 19:72:@5332.4]
  wire [7:0] _T_6845; // @[Mux.scala 19:72:@5333.4]
  wire [7:0] _T_6846; // @[Mux.scala 19:72:@5334.4]
  wire [7:0] _T_7088; // @[Mux.scala 19:72:@5452.4]
  wire [7:0] _T_7090; // @[Mux.scala 19:72:@5453.4]
  wire [7:0] _T_7097; // @[Mux.scala 19:72:@5460.4]
  wire [7:0] _T_7099; // @[Mux.scala 19:72:@5461.4]
  wire [7:0] _T_7106; // @[Mux.scala 19:72:@5468.4]
  wire [7:0] _T_7108; // @[Mux.scala 19:72:@5469.4]
  wire [7:0] _T_7115; // @[Mux.scala 19:72:@5476.4]
  wire [7:0] _T_7117; // @[Mux.scala 19:72:@5477.4]
  wire [7:0] _T_7124; // @[Mux.scala 19:72:@5484.4]
  wire [7:0] _T_7126; // @[Mux.scala 19:72:@5485.4]
  wire [7:0] _T_7133; // @[Mux.scala 19:72:@5492.4]
  wire [7:0] _T_7135; // @[Mux.scala 19:72:@5493.4]
  wire [7:0] _T_7142; // @[Mux.scala 19:72:@5500.4]
  wire [7:0] _T_7144; // @[Mux.scala 19:72:@5501.4]
  wire [7:0] _T_7151; // @[Mux.scala 19:72:@5508.4]
  wire [7:0] _T_7153; // @[Mux.scala 19:72:@5509.4]
  wire [7:0] _T_7154; // @[Mux.scala 19:72:@5510.4]
  wire [7:0] _T_7155; // @[Mux.scala 19:72:@5511.4]
  wire [7:0] _T_7156; // @[Mux.scala 19:72:@5512.4]
  wire [7:0] _T_7157; // @[Mux.scala 19:72:@5513.4]
  wire [7:0] _T_7158; // @[Mux.scala 19:72:@5514.4]
  wire [7:0] _T_7159; // @[Mux.scala 19:72:@5515.4]
  wire [7:0] _T_7160; // @[Mux.scala 19:72:@5516.4]
  wire [7:0] _T_7402; // @[Mux.scala 19:72:@5634.4]
  wire [7:0] _T_7404; // @[Mux.scala 19:72:@5635.4]
  wire [7:0] _T_7411; // @[Mux.scala 19:72:@5642.4]
  wire [7:0] _T_7413; // @[Mux.scala 19:72:@5643.4]
  wire [7:0] _T_7420; // @[Mux.scala 19:72:@5650.4]
  wire [7:0] _T_7422; // @[Mux.scala 19:72:@5651.4]
  wire [7:0] _T_7429; // @[Mux.scala 19:72:@5658.4]
  wire [7:0] _T_7431; // @[Mux.scala 19:72:@5659.4]
  wire [7:0] _T_7438; // @[Mux.scala 19:72:@5666.4]
  wire [7:0] _T_7440; // @[Mux.scala 19:72:@5667.4]
  wire [7:0] _T_7447; // @[Mux.scala 19:72:@5674.4]
  wire [7:0] _T_7449; // @[Mux.scala 19:72:@5675.4]
  wire [7:0] _T_7456; // @[Mux.scala 19:72:@5682.4]
  wire [7:0] _T_7458; // @[Mux.scala 19:72:@5683.4]
  wire [7:0] _T_7465; // @[Mux.scala 19:72:@5690.4]
  wire [7:0] _T_7467; // @[Mux.scala 19:72:@5691.4]
  wire [7:0] _T_7468; // @[Mux.scala 19:72:@5692.4]
  wire [7:0] _T_7469; // @[Mux.scala 19:72:@5693.4]
  wire [7:0] _T_7470; // @[Mux.scala 19:72:@5694.4]
  wire [7:0] _T_7471; // @[Mux.scala 19:72:@5695.4]
  wire [7:0] _T_7472; // @[Mux.scala 19:72:@5696.4]
  wire [7:0] _T_7473; // @[Mux.scala 19:72:@5697.4]
  wire [7:0] _T_7474; // @[Mux.scala 19:72:@5698.4]
  wire [7:0] _T_7716; // @[Mux.scala 19:72:@5816.4]
  wire [7:0] _T_7718; // @[Mux.scala 19:72:@5817.4]
  wire [7:0] _T_7725; // @[Mux.scala 19:72:@5824.4]
  wire [7:0] _T_7727; // @[Mux.scala 19:72:@5825.4]
  wire [7:0] _T_7734; // @[Mux.scala 19:72:@5832.4]
  wire [7:0] _T_7736; // @[Mux.scala 19:72:@5833.4]
  wire [7:0] _T_7743; // @[Mux.scala 19:72:@5840.4]
  wire [7:0] _T_7745; // @[Mux.scala 19:72:@5841.4]
  wire [7:0] _T_7752; // @[Mux.scala 19:72:@5848.4]
  wire [7:0] _T_7754; // @[Mux.scala 19:72:@5849.4]
  wire [7:0] _T_7761; // @[Mux.scala 19:72:@5856.4]
  wire [7:0] _T_7763; // @[Mux.scala 19:72:@5857.4]
  wire [7:0] _T_7770; // @[Mux.scala 19:72:@5864.4]
  wire [7:0] _T_7772; // @[Mux.scala 19:72:@5865.4]
  wire [7:0] _T_7779; // @[Mux.scala 19:72:@5872.4]
  wire [7:0] _T_7781; // @[Mux.scala 19:72:@5873.4]
  wire [7:0] _T_7782; // @[Mux.scala 19:72:@5874.4]
  wire [7:0] _T_7783; // @[Mux.scala 19:72:@5875.4]
  wire [7:0] _T_7784; // @[Mux.scala 19:72:@5876.4]
  wire [7:0] _T_7785; // @[Mux.scala 19:72:@5877.4]
  wire [7:0] _T_7786; // @[Mux.scala 19:72:@5878.4]
  wire [7:0] _T_7787; // @[Mux.scala 19:72:@5879.4]
  wire [7:0] _T_7788; // @[Mux.scala 19:72:@5880.4]
  wire [7:0] _T_8030; // @[Mux.scala 19:72:@5998.4]
  wire [7:0] _T_8032; // @[Mux.scala 19:72:@5999.4]
  wire [7:0] _T_8039; // @[Mux.scala 19:72:@6006.4]
  wire [7:0] _T_8041; // @[Mux.scala 19:72:@6007.4]
  wire [7:0] _T_8048; // @[Mux.scala 19:72:@6014.4]
  wire [7:0] _T_8050; // @[Mux.scala 19:72:@6015.4]
  wire [7:0] _T_8057; // @[Mux.scala 19:72:@6022.4]
  wire [7:0] _T_8059; // @[Mux.scala 19:72:@6023.4]
  wire [7:0] _T_8066; // @[Mux.scala 19:72:@6030.4]
  wire [7:0] _T_8068; // @[Mux.scala 19:72:@6031.4]
  wire [7:0] _T_8075; // @[Mux.scala 19:72:@6038.4]
  wire [7:0] _T_8077; // @[Mux.scala 19:72:@6039.4]
  wire [7:0] _T_8084; // @[Mux.scala 19:72:@6046.4]
  wire [7:0] _T_8086; // @[Mux.scala 19:72:@6047.4]
  wire [7:0] _T_8093; // @[Mux.scala 19:72:@6054.4]
  wire [7:0] _T_8095; // @[Mux.scala 19:72:@6055.4]
  wire [7:0] _T_8096; // @[Mux.scala 19:72:@6056.4]
  wire [7:0] _T_8097; // @[Mux.scala 19:72:@6057.4]
  wire [7:0] _T_8098; // @[Mux.scala 19:72:@6058.4]
  wire [7:0] _T_8099; // @[Mux.scala 19:72:@6059.4]
  wire [7:0] _T_8100; // @[Mux.scala 19:72:@6060.4]
  wire [7:0] _T_8101; // @[Mux.scala 19:72:@6061.4]
  wire [7:0] _T_8102; // @[Mux.scala 19:72:@6062.4]
  wire [7:0] _T_8344; // @[Mux.scala 19:72:@6180.4]
  wire [7:0] _T_8346; // @[Mux.scala 19:72:@6181.4]
  wire [7:0] _T_8353; // @[Mux.scala 19:72:@6188.4]
  wire [7:0] _T_8355; // @[Mux.scala 19:72:@6189.4]
  wire [7:0] _T_8362; // @[Mux.scala 19:72:@6196.4]
  wire [7:0] _T_8364; // @[Mux.scala 19:72:@6197.4]
  wire [7:0] _T_8371; // @[Mux.scala 19:72:@6204.4]
  wire [7:0] _T_8373; // @[Mux.scala 19:72:@6205.4]
  wire [7:0] _T_8380; // @[Mux.scala 19:72:@6212.4]
  wire [7:0] _T_8382; // @[Mux.scala 19:72:@6213.4]
  wire [7:0] _T_8389; // @[Mux.scala 19:72:@6220.4]
  wire [7:0] _T_8391; // @[Mux.scala 19:72:@6221.4]
  wire [7:0] _T_8398; // @[Mux.scala 19:72:@6228.4]
  wire [7:0] _T_8400; // @[Mux.scala 19:72:@6229.4]
  wire [7:0] _T_8407; // @[Mux.scala 19:72:@6236.4]
  wire [7:0] _T_8409; // @[Mux.scala 19:72:@6237.4]
  wire [7:0] _T_8410; // @[Mux.scala 19:72:@6238.4]
  wire [7:0] _T_8411; // @[Mux.scala 19:72:@6239.4]
  wire [7:0] _T_8412; // @[Mux.scala 19:72:@6240.4]
  wire [7:0] _T_8413; // @[Mux.scala 19:72:@6241.4]
  wire [7:0] _T_8414; // @[Mux.scala 19:72:@6242.4]
  wire [7:0] _T_8415; // @[Mux.scala 19:72:@6243.4]
  wire [7:0] _T_8416; // @[Mux.scala 19:72:@6244.4]
  reg  conflictPReg_0_0; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_83;
  reg  conflictPReg_0_1; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_84;
  reg  conflictPReg_0_2; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_85;
  reg  conflictPReg_0_3; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_86;
  reg  conflictPReg_0_4; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_87;
  reg  conflictPReg_0_5; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_88;
  reg  conflictPReg_0_6; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_89;
  reg  conflictPReg_0_7; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_90;
  reg  conflictPReg_1_0; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_91;
  reg  conflictPReg_1_1; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_92;
  reg  conflictPReg_1_2; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_93;
  reg  conflictPReg_1_3; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_94;
  reg  conflictPReg_1_4; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_95;
  reg  conflictPReg_1_5; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_96;
  reg  conflictPReg_1_6; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_97;
  reg  conflictPReg_1_7; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_98;
  reg  conflictPReg_2_0; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_99;
  reg  conflictPReg_2_1; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_100;
  reg  conflictPReg_2_2; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_101;
  reg  conflictPReg_2_3; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_102;
  reg  conflictPReg_2_4; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_103;
  reg  conflictPReg_2_5; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_104;
  reg  conflictPReg_2_6; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_105;
  reg  conflictPReg_2_7; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_106;
  reg  conflictPReg_3_0; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_107;
  reg  conflictPReg_3_1; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_108;
  reg  conflictPReg_3_2; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_109;
  reg  conflictPReg_3_3; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_110;
  reg  conflictPReg_3_4; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_111;
  reg  conflictPReg_3_5; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_112;
  reg  conflictPReg_3_6; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_113;
  reg  conflictPReg_3_7; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_114;
  reg  conflictPReg_4_0; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_115;
  reg  conflictPReg_4_1; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_116;
  reg  conflictPReg_4_2; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_117;
  reg  conflictPReg_4_3; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_118;
  reg  conflictPReg_4_4; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_119;
  reg  conflictPReg_4_5; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_120;
  reg  conflictPReg_4_6; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_121;
  reg  conflictPReg_4_7; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_122;
  reg  conflictPReg_5_0; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_123;
  reg  conflictPReg_5_1; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_124;
  reg  conflictPReg_5_2; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_125;
  reg  conflictPReg_5_3; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_126;
  reg  conflictPReg_5_4; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_127;
  reg  conflictPReg_5_5; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_128;
  reg  conflictPReg_5_6; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_129;
  reg  conflictPReg_5_7; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_130;
  reg  conflictPReg_6_0; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_131;
  reg  conflictPReg_6_1; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_132;
  reg  conflictPReg_6_2; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_133;
  reg  conflictPReg_6_3; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_134;
  reg  conflictPReg_6_4; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_135;
  reg  conflictPReg_6_5; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_136;
  reg  conflictPReg_6_6; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_137;
  reg  conflictPReg_6_7; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_138;
  reg  conflictPReg_7_0; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_139;
  reg  conflictPReg_7_1; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_140;
  reg  conflictPReg_7_2; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_141;
  reg  conflictPReg_7_3; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_142;
  reg  conflictPReg_7_4; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_143;
  reg  conflictPReg_7_5; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_144;
  reg  conflictPReg_7_6; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_145;
  reg  conflictPReg_7_7; // @[LoadQueue.scala 166:29:@6329.4]
  reg [31:0] _RAND_146;
  wire [7:0] _T_14526; // @[Mux.scala 19:72:@6492.4]
  wire [7:0] _T_14528; // @[Mux.scala 19:72:@6493.4]
  wire [7:0] _T_14535; // @[Mux.scala 19:72:@6500.4]
  wire [7:0] _T_14537; // @[Mux.scala 19:72:@6501.4]
  wire [7:0] _T_14544; // @[Mux.scala 19:72:@6508.4]
  wire [7:0] _T_14546; // @[Mux.scala 19:72:@6509.4]
  wire [7:0] _T_14553; // @[Mux.scala 19:72:@6516.4]
  wire [7:0] _T_14555; // @[Mux.scala 19:72:@6517.4]
  wire [7:0] _T_14562; // @[Mux.scala 19:72:@6524.4]
  wire [7:0] _T_14564; // @[Mux.scala 19:72:@6525.4]
  wire [7:0] _T_14571; // @[Mux.scala 19:72:@6532.4]
  wire [7:0] _T_14573; // @[Mux.scala 19:72:@6533.4]
  wire [7:0] _T_14580; // @[Mux.scala 19:72:@6540.4]
  wire [7:0] _T_14582; // @[Mux.scala 19:72:@6541.4]
  wire [7:0] _T_14589; // @[Mux.scala 19:72:@6548.4]
  wire [7:0] _T_14591; // @[Mux.scala 19:72:@6549.4]
  wire [7:0] _T_14592; // @[Mux.scala 19:72:@6550.4]
  wire [7:0] _T_14593; // @[Mux.scala 19:72:@6551.4]
  wire [7:0] _T_14594; // @[Mux.scala 19:72:@6552.4]
  wire [7:0] _T_14595; // @[Mux.scala 19:72:@6553.4]
  wire [7:0] _T_14596; // @[Mux.scala 19:72:@6554.4]
  wire [7:0] _T_14597; // @[Mux.scala 19:72:@6555.4]
  wire [7:0] _T_14598; // @[Mux.scala 19:72:@6556.4]
  wire [7:0] _T_14840; // @[Mux.scala 19:72:@6674.4]
  wire [7:0] _T_14842; // @[Mux.scala 19:72:@6675.4]
  wire [7:0] _T_14849; // @[Mux.scala 19:72:@6682.4]
  wire [7:0] _T_14851; // @[Mux.scala 19:72:@6683.4]
  wire [7:0] _T_14858; // @[Mux.scala 19:72:@6690.4]
  wire [7:0] _T_14860; // @[Mux.scala 19:72:@6691.4]
  wire [7:0] _T_14867; // @[Mux.scala 19:72:@6698.4]
  wire [7:0] _T_14869; // @[Mux.scala 19:72:@6699.4]
  wire [7:0] _T_14876; // @[Mux.scala 19:72:@6706.4]
  wire [7:0] _T_14878; // @[Mux.scala 19:72:@6707.4]
  wire [7:0] _T_14885; // @[Mux.scala 19:72:@6714.4]
  wire [7:0] _T_14887; // @[Mux.scala 19:72:@6715.4]
  wire [7:0] _T_14894; // @[Mux.scala 19:72:@6722.4]
  wire [7:0] _T_14896; // @[Mux.scala 19:72:@6723.4]
  wire [7:0] _T_14903; // @[Mux.scala 19:72:@6730.4]
  wire [7:0] _T_14905; // @[Mux.scala 19:72:@6731.4]
  wire [7:0] _T_14906; // @[Mux.scala 19:72:@6732.4]
  wire [7:0] _T_14907; // @[Mux.scala 19:72:@6733.4]
  wire [7:0] _T_14908; // @[Mux.scala 19:72:@6734.4]
  wire [7:0] _T_14909; // @[Mux.scala 19:72:@6735.4]
  wire [7:0] _T_14910; // @[Mux.scala 19:72:@6736.4]
  wire [7:0] _T_14911; // @[Mux.scala 19:72:@6737.4]
  wire [7:0] _T_14912; // @[Mux.scala 19:72:@6738.4]
  wire [7:0] _T_15154; // @[Mux.scala 19:72:@6856.4]
  wire [7:0] _T_15156; // @[Mux.scala 19:72:@6857.4]
  wire [7:0] _T_15163; // @[Mux.scala 19:72:@6864.4]
  wire [7:0] _T_15165; // @[Mux.scala 19:72:@6865.4]
  wire [7:0] _T_15172; // @[Mux.scala 19:72:@6872.4]
  wire [7:0] _T_15174; // @[Mux.scala 19:72:@6873.4]
  wire [7:0] _T_15181; // @[Mux.scala 19:72:@6880.4]
  wire [7:0] _T_15183; // @[Mux.scala 19:72:@6881.4]
  wire [7:0] _T_15190; // @[Mux.scala 19:72:@6888.4]
  wire [7:0] _T_15192; // @[Mux.scala 19:72:@6889.4]
  wire [7:0] _T_15199; // @[Mux.scala 19:72:@6896.4]
  wire [7:0] _T_15201; // @[Mux.scala 19:72:@6897.4]
  wire [7:0] _T_15208; // @[Mux.scala 19:72:@6904.4]
  wire [7:0] _T_15210; // @[Mux.scala 19:72:@6905.4]
  wire [7:0] _T_15217; // @[Mux.scala 19:72:@6912.4]
  wire [7:0] _T_15219; // @[Mux.scala 19:72:@6913.4]
  wire [7:0] _T_15220; // @[Mux.scala 19:72:@6914.4]
  wire [7:0] _T_15221; // @[Mux.scala 19:72:@6915.4]
  wire [7:0] _T_15222; // @[Mux.scala 19:72:@6916.4]
  wire [7:0] _T_15223; // @[Mux.scala 19:72:@6917.4]
  wire [7:0] _T_15224; // @[Mux.scala 19:72:@6918.4]
  wire [7:0] _T_15225; // @[Mux.scala 19:72:@6919.4]
  wire [7:0] _T_15226; // @[Mux.scala 19:72:@6920.4]
  wire [7:0] _T_15468; // @[Mux.scala 19:72:@7038.4]
  wire [7:0] _T_15470; // @[Mux.scala 19:72:@7039.4]
  wire [7:0] _T_15477; // @[Mux.scala 19:72:@7046.4]
  wire [7:0] _T_15479; // @[Mux.scala 19:72:@7047.4]
  wire [7:0] _T_15486; // @[Mux.scala 19:72:@7054.4]
  wire [7:0] _T_15488; // @[Mux.scala 19:72:@7055.4]
  wire [7:0] _T_15495; // @[Mux.scala 19:72:@7062.4]
  wire [7:0] _T_15497; // @[Mux.scala 19:72:@7063.4]
  wire [7:0] _T_15504; // @[Mux.scala 19:72:@7070.4]
  wire [7:0] _T_15506; // @[Mux.scala 19:72:@7071.4]
  wire [7:0] _T_15513; // @[Mux.scala 19:72:@7078.4]
  wire [7:0] _T_15515; // @[Mux.scala 19:72:@7079.4]
  wire [7:0] _T_15522; // @[Mux.scala 19:72:@7086.4]
  wire [7:0] _T_15524; // @[Mux.scala 19:72:@7087.4]
  wire [7:0] _T_15531; // @[Mux.scala 19:72:@7094.4]
  wire [7:0] _T_15533; // @[Mux.scala 19:72:@7095.4]
  wire [7:0] _T_15534; // @[Mux.scala 19:72:@7096.4]
  wire [7:0] _T_15535; // @[Mux.scala 19:72:@7097.4]
  wire [7:0] _T_15536; // @[Mux.scala 19:72:@7098.4]
  wire [7:0] _T_15537; // @[Mux.scala 19:72:@7099.4]
  wire [7:0] _T_15538; // @[Mux.scala 19:72:@7100.4]
  wire [7:0] _T_15539; // @[Mux.scala 19:72:@7101.4]
  wire [7:0] _T_15540; // @[Mux.scala 19:72:@7102.4]
  wire [7:0] _T_15782; // @[Mux.scala 19:72:@7220.4]
  wire [7:0] _T_15784; // @[Mux.scala 19:72:@7221.4]
  wire [7:0] _T_15791; // @[Mux.scala 19:72:@7228.4]
  wire [7:0] _T_15793; // @[Mux.scala 19:72:@7229.4]
  wire [7:0] _T_15800; // @[Mux.scala 19:72:@7236.4]
  wire [7:0] _T_15802; // @[Mux.scala 19:72:@7237.4]
  wire [7:0] _T_15809; // @[Mux.scala 19:72:@7244.4]
  wire [7:0] _T_15811; // @[Mux.scala 19:72:@7245.4]
  wire [7:0] _T_15818; // @[Mux.scala 19:72:@7252.4]
  wire [7:0] _T_15820; // @[Mux.scala 19:72:@7253.4]
  wire [7:0] _T_15827; // @[Mux.scala 19:72:@7260.4]
  wire [7:0] _T_15829; // @[Mux.scala 19:72:@7261.4]
  wire [7:0] _T_15836; // @[Mux.scala 19:72:@7268.4]
  wire [7:0] _T_15838; // @[Mux.scala 19:72:@7269.4]
  wire [7:0] _T_15845; // @[Mux.scala 19:72:@7276.4]
  wire [7:0] _T_15847; // @[Mux.scala 19:72:@7277.4]
  wire [7:0] _T_15848; // @[Mux.scala 19:72:@7278.4]
  wire [7:0] _T_15849; // @[Mux.scala 19:72:@7279.4]
  wire [7:0] _T_15850; // @[Mux.scala 19:72:@7280.4]
  wire [7:0] _T_15851; // @[Mux.scala 19:72:@7281.4]
  wire [7:0] _T_15852; // @[Mux.scala 19:72:@7282.4]
  wire [7:0] _T_15853; // @[Mux.scala 19:72:@7283.4]
  wire [7:0] _T_15854; // @[Mux.scala 19:72:@7284.4]
  wire [7:0] _T_16096; // @[Mux.scala 19:72:@7402.4]
  wire [7:0] _T_16098; // @[Mux.scala 19:72:@7403.4]
  wire [7:0] _T_16105; // @[Mux.scala 19:72:@7410.4]
  wire [7:0] _T_16107; // @[Mux.scala 19:72:@7411.4]
  wire [7:0] _T_16114; // @[Mux.scala 19:72:@7418.4]
  wire [7:0] _T_16116; // @[Mux.scala 19:72:@7419.4]
  wire [7:0] _T_16123; // @[Mux.scala 19:72:@7426.4]
  wire [7:0] _T_16125; // @[Mux.scala 19:72:@7427.4]
  wire [7:0] _T_16132; // @[Mux.scala 19:72:@7434.4]
  wire [7:0] _T_16134; // @[Mux.scala 19:72:@7435.4]
  wire [7:0] _T_16141; // @[Mux.scala 19:72:@7442.4]
  wire [7:0] _T_16143; // @[Mux.scala 19:72:@7443.4]
  wire [7:0] _T_16150; // @[Mux.scala 19:72:@7450.4]
  wire [7:0] _T_16152; // @[Mux.scala 19:72:@7451.4]
  wire [7:0] _T_16159; // @[Mux.scala 19:72:@7458.4]
  wire [7:0] _T_16161; // @[Mux.scala 19:72:@7459.4]
  wire [7:0] _T_16162; // @[Mux.scala 19:72:@7460.4]
  wire [7:0] _T_16163; // @[Mux.scala 19:72:@7461.4]
  wire [7:0] _T_16164; // @[Mux.scala 19:72:@7462.4]
  wire [7:0] _T_16165; // @[Mux.scala 19:72:@7463.4]
  wire [7:0] _T_16166; // @[Mux.scala 19:72:@7464.4]
  wire [7:0] _T_16167; // @[Mux.scala 19:72:@7465.4]
  wire [7:0] _T_16168; // @[Mux.scala 19:72:@7466.4]
  wire [7:0] _T_16410; // @[Mux.scala 19:72:@7584.4]
  wire [7:0] _T_16412; // @[Mux.scala 19:72:@7585.4]
  wire [7:0] _T_16419; // @[Mux.scala 19:72:@7592.4]
  wire [7:0] _T_16421; // @[Mux.scala 19:72:@7593.4]
  wire [7:0] _T_16428; // @[Mux.scala 19:72:@7600.4]
  wire [7:0] _T_16430; // @[Mux.scala 19:72:@7601.4]
  wire [7:0] _T_16437; // @[Mux.scala 19:72:@7608.4]
  wire [7:0] _T_16439; // @[Mux.scala 19:72:@7609.4]
  wire [7:0] _T_16446; // @[Mux.scala 19:72:@7616.4]
  wire [7:0] _T_16448; // @[Mux.scala 19:72:@7617.4]
  wire [7:0] _T_16455; // @[Mux.scala 19:72:@7624.4]
  wire [7:0] _T_16457; // @[Mux.scala 19:72:@7625.4]
  wire [7:0] _T_16464; // @[Mux.scala 19:72:@7632.4]
  wire [7:0] _T_16466; // @[Mux.scala 19:72:@7633.4]
  wire [7:0] _T_16473; // @[Mux.scala 19:72:@7640.4]
  wire [7:0] _T_16475; // @[Mux.scala 19:72:@7641.4]
  wire [7:0] _T_16476; // @[Mux.scala 19:72:@7642.4]
  wire [7:0] _T_16477; // @[Mux.scala 19:72:@7643.4]
  wire [7:0] _T_16478; // @[Mux.scala 19:72:@7644.4]
  wire [7:0] _T_16479; // @[Mux.scala 19:72:@7645.4]
  wire [7:0] _T_16480; // @[Mux.scala 19:72:@7646.4]
  wire [7:0] _T_16481; // @[Mux.scala 19:72:@7647.4]
  wire [7:0] _T_16482; // @[Mux.scala 19:72:@7648.4]
  wire [7:0] _T_16724; // @[Mux.scala 19:72:@7766.4]
  wire [7:0] _T_16726; // @[Mux.scala 19:72:@7767.4]
  wire [7:0] _T_16733; // @[Mux.scala 19:72:@7774.4]
  wire [7:0] _T_16735; // @[Mux.scala 19:72:@7775.4]
  wire [7:0] _T_16742; // @[Mux.scala 19:72:@7782.4]
  wire [7:0] _T_16744; // @[Mux.scala 19:72:@7783.4]
  wire [7:0] _T_16751; // @[Mux.scala 19:72:@7790.4]
  wire [7:0] _T_16753; // @[Mux.scala 19:72:@7791.4]
  wire [7:0] _T_16760; // @[Mux.scala 19:72:@7798.4]
  wire [7:0] _T_16762; // @[Mux.scala 19:72:@7799.4]
  wire [7:0] _T_16769; // @[Mux.scala 19:72:@7806.4]
  wire [7:0] _T_16771; // @[Mux.scala 19:72:@7807.4]
  wire [7:0] _T_16778; // @[Mux.scala 19:72:@7814.4]
  wire [7:0] _T_16780; // @[Mux.scala 19:72:@7815.4]
  wire [7:0] _T_16787; // @[Mux.scala 19:72:@7822.4]
  wire [7:0] _T_16789; // @[Mux.scala 19:72:@7823.4]
  wire [7:0] _T_16790; // @[Mux.scala 19:72:@7824.4]
  wire [7:0] _T_16791; // @[Mux.scala 19:72:@7825.4]
  wire [7:0] _T_16792; // @[Mux.scala 19:72:@7826.4]
  wire [7:0] _T_16793; // @[Mux.scala 19:72:@7827.4]
  wire [7:0] _T_16794; // @[Mux.scala 19:72:@7828.4]
  wire [7:0] _T_16795; // @[Mux.scala 19:72:@7829.4]
  wire [7:0] _T_16796; // @[Mux.scala 19:72:@7830.4]
  reg  storeAddrNotKnownFlagsPReg_0_0; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_147;
  reg  storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_148;
  reg  storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_149;
  reg  storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_150;
  reg  storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_151;
  reg  storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_152;
  reg  storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_153;
  reg  storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_154;
  reg  storeAddrNotKnownFlagsPReg_1_0; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_155;
  reg  storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_156;
  reg  storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_157;
  reg  storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_158;
  reg  storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_159;
  reg  storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_160;
  reg  storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_161;
  reg  storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_162;
  reg  storeAddrNotKnownFlagsPReg_2_0; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_163;
  reg  storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_164;
  reg  storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_165;
  reg  storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_166;
  reg  storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_167;
  reg  storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_168;
  reg  storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_169;
  reg  storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_170;
  reg  storeAddrNotKnownFlagsPReg_3_0; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_171;
  reg  storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_172;
  reg  storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_173;
  reg  storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_174;
  reg  storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_175;
  reg  storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_176;
  reg  storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_177;
  reg  storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_178;
  reg  storeAddrNotKnownFlagsPReg_4_0; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_179;
  reg  storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_180;
  reg  storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_181;
  reg  storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_182;
  reg  storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_183;
  reg  storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_184;
  reg  storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_185;
  reg  storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_186;
  reg  storeAddrNotKnownFlagsPReg_5_0; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_187;
  reg  storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_188;
  reg  storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_189;
  reg  storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_190;
  reg  storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_191;
  reg  storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_192;
  reg  storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_193;
  reg  storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_194;
  reg  storeAddrNotKnownFlagsPReg_6_0; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_195;
  reg  storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_196;
  reg  storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_197;
  reg  storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_198;
  reg  storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_199;
  reg  storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_200;
  reg  storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_201;
  reg  storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_202;
  reg  storeAddrNotKnownFlagsPReg_7_0; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_203;
  reg  storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_204;
  reg  storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_205;
  reg  storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_206;
  reg  storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_207;
  reg  storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_208;
  reg  storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_209;
  reg  storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 167:43:@7915.4]
  reg [31:0] _RAND_210;
  reg  shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 168:42:@7980.4]
  reg [31:0] _RAND_211;
  reg  shiftedStoreDataKnownPReg_1; // @[LoadQueue.scala 168:42:@7980.4]
  reg [31:0] _RAND_212;
  reg  shiftedStoreDataKnownPReg_2; // @[LoadQueue.scala 168:42:@7980.4]
  reg [31:0] _RAND_213;
  reg  shiftedStoreDataKnownPReg_3; // @[LoadQueue.scala 168:42:@7980.4]
  reg [31:0] _RAND_214;
  reg  shiftedStoreDataKnownPReg_4; // @[LoadQueue.scala 168:42:@7980.4]
  reg [31:0] _RAND_215;
  reg  shiftedStoreDataKnownPReg_5; // @[LoadQueue.scala 168:42:@7980.4]
  reg [31:0] _RAND_216;
  reg  shiftedStoreDataKnownPReg_6; // @[LoadQueue.scala 168:42:@7980.4]
  reg [31:0] _RAND_217;
  reg  shiftedStoreDataKnownPReg_7; // @[LoadQueue.scala 168:42:@7980.4]
  reg [31:0] _RAND_218;
  reg [31:0] shiftedStoreDataQPreg_0; // @[LoadQueue.scala 169:38:@7989.4]
  reg [31:0] _RAND_219;
  reg [31:0] shiftedStoreDataQPreg_1; // @[LoadQueue.scala 169:38:@7989.4]
  reg [31:0] _RAND_220;
  reg [31:0] shiftedStoreDataQPreg_2; // @[LoadQueue.scala 169:38:@7989.4]
  reg [31:0] _RAND_221;
  reg [31:0] shiftedStoreDataQPreg_3; // @[LoadQueue.scala 169:38:@7989.4]
  reg [31:0] _RAND_222;
  reg [31:0] shiftedStoreDataQPreg_4; // @[LoadQueue.scala 169:38:@7989.4]
  reg [31:0] _RAND_223;
  reg [31:0] shiftedStoreDataQPreg_5; // @[LoadQueue.scala 169:38:@7989.4]
  reg [31:0] _RAND_224;
  reg [31:0] shiftedStoreDataQPreg_6; // @[LoadQueue.scala 169:38:@7989.4]
  reg [31:0] _RAND_225;
  reg [31:0] shiftedStoreDataQPreg_7; // @[LoadQueue.scala 169:38:@7989.4]
  reg [31:0] _RAND_226;
  reg  addrKnownPReg_0; // @[LoadQueue.scala 170:30:@7998.4]
  reg [31:0] _RAND_227;
  reg  addrKnownPReg_1; // @[LoadQueue.scala 170:30:@7998.4]
  reg [31:0] _RAND_228;
  reg  addrKnownPReg_2; // @[LoadQueue.scala 170:30:@7998.4]
  reg [31:0] _RAND_229;
  reg  addrKnownPReg_3; // @[LoadQueue.scala 170:30:@7998.4]
  reg [31:0] _RAND_230;
  reg  addrKnownPReg_4; // @[LoadQueue.scala 170:30:@7998.4]
  reg [31:0] _RAND_231;
  reg  addrKnownPReg_5; // @[LoadQueue.scala 170:30:@7998.4]
  reg [31:0] _RAND_232;
  reg  addrKnownPReg_6; // @[LoadQueue.scala 170:30:@7998.4]
  reg [31:0] _RAND_233;
  reg  addrKnownPReg_7; // @[LoadQueue.scala 170:30:@7998.4]
  reg [31:0] _RAND_234;
  reg  dataKnownPReg_0; // @[LoadQueue.scala 171:30:@8007.4]
  reg [31:0] _RAND_235;
  reg  dataKnownPReg_1; // @[LoadQueue.scala 171:30:@8007.4]
  reg [31:0] _RAND_236;
  reg  dataKnownPReg_2; // @[LoadQueue.scala 171:30:@8007.4]
  reg [31:0] _RAND_237;
  reg  dataKnownPReg_3; // @[LoadQueue.scala 171:30:@8007.4]
  reg [31:0] _RAND_238;
  reg  dataKnownPReg_4; // @[LoadQueue.scala 171:30:@8007.4]
  reg [31:0] _RAND_239;
  reg  dataKnownPReg_5; // @[LoadQueue.scala 171:30:@8007.4]
  reg [31:0] _RAND_240;
  reg  dataKnownPReg_6; // @[LoadQueue.scala 171:30:@8007.4]
  reg [31:0] _RAND_241;
  reg  dataKnownPReg_7; // @[LoadQueue.scala 171:30:@8007.4]
  reg [31:0] _RAND_242;
  wire [1:0] _T_23556; // @[LoadQueue.scala 191:60:@8047.4]
  wire [1:0] _T_23557; // @[LoadQueue.scala 191:60:@8048.4]
  wire [2:0] _T_23558; // @[LoadQueue.scala 191:60:@8049.4]
  wire [2:0] _T_23559; // @[LoadQueue.scala 191:60:@8050.4]
  wire [2:0] _T_23560; // @[LoadQueue.scala 191:60:@8051.4]
  wire [2:0] _T_23561; // @[LoadQueue.scala 191:60:@8052.4]
  wire  _T_23564; // @[LoadQueue.scala 192:43:@8054.4]
  wire  _T_23565; // @[LoadQueue.scala 192:43:@8055.4]
  wire  _T_23566; // @[LoadQueue.scala 192:43:@8056.4]
  wire  _T_23567; // @[LoadQueue.scala 192:43:@8057.4]
  wire  _T_23568; // @[LoadQueue.scala 192:43:@8058.4]
  wire  _T_23569; // @[LoadQueue.scala 192:43:@8059.4]
  wire  _T_23570; // @[LoadQueue.scala 192:43:@8060.4]
  wire  _GEN_240; // @[LoadQueue.scala 193:43:@8062.6]
  wire  _GEN_241; // @[LoadQueue.scala 193:43:@8062.6]
  wire  _GEN_242; // @[LoadQueue.scala 193:43:@8062.6]
  wire  _GEN_243; // @[LoadQueue.scala 193:43:@8062.6]
  wire  _GEN_244; // @[LoadQueue.scala 193:43:@8062.6]
  wire  _GEN_245; // @[LoadQueue.scala 193:43:@8062.6]
  wire  _GEN_246; // @[LoadQueue.scala 193:43:@8062.6]
  wire  _GEN_247; // @[LoadQueue.scala 193:43:@8062.6]
  wire  _GEN_249; // @[LoadQueue.scala 194:31:@8063.6]
  wire  _GEN_250; // @[LoadQueue.scala 194:31:@8063.6]
  wire  _GEN_251; // @[LoadQueue.scala 194:31:@8063.6]
  wire  _GEN_252; // @[LoadQueue.scala 194:31:@8063.6]
  wire  _GEN_253; // @[LoadQueue.scala 194:31:@8063.6]
  wire  _GEN_254; // @[LoadQueue.scala 194:31:@8063.6]
  wire  _GEN_255; // @[LoadQueue.scala 194:31:@8063.6]
  wire [31:0] _GEN_257; // @[LoadQueue.scala 195:31:@8064.6]
  wire [31:0] _GEN_258; // @[LoadQueue.scala 195:31:@8064.6]
  wire [31:0] _GEN_259; // @[LoadQueue.scala 195:31:@8064.6]
  wire [31:0] _GEN_260; // @[LoadQueue.scala 195:31:@8064.6]
  wire [31:0] _GEN_261; // @[LoadQueue.scala 195:31:@8064.6]
  wire [31:0] _GEN_262; // @[LoadQueue.scala 195:31:@8064.6]
  wire [31:0] _GEN_263; // @[LoadQueue.scala 195:31:@8064.6]
  wire  lastConflict_0_0; // @[LoadQueue.scala 192:53:@8061.4]
  wire  lastConflict_0_1; // @[LoadQueue.scala 192:53:@8061.4]
  wire  lastConflict_0_2; // @[LoadQueue.scala 192:53:@8061.4]
  wire  lastConflict_0_3; // @[LoadQueue.scala 192:53:@8061.4]
  wire  lastConflict_0_4; // @[LoadQueue.scala 192:53:@8061.4]
  wire  lastConflict_0_5; // @[LoadQueue.scala 192:53:@8061.4]
  wire  lastConflict_0_6; // @[LoadQueue.scala 192:53:@8061.4]
  wire  lastConflict_0_7; // @[LoadQueue.scala 192:53:@8061.4]
  wire  canBypass_0; // @[LoadQueue.scala 192:53:@8061.4]
  wire [31:0] bypassVal_0; // @[LoadQueue.scala 192:53:@8061.4]
  wire [1:0] _T_23636; // @[LoadQueue.scala 191:60:@8094.4]
  wire [1:0] _T_23637; // @[LoadQueue.scala 191:60:@8095.4]
  wire [2:0] _T_23638; // @[LoadQueue.scala 191:60:@8096.4]
  wire [2:0] _T_23639; // @[LoadQueue.scala 191:60:@8097.4]
  wire [2:0] _T_23640; // @[LoadQueue.scala 191:60:@8098.4]
  wire [2:0] _T_23641; // @[LoadQueue.scala 191:60:@8099.4]
  wire  _T_23644; // @[LoadQueue.scala 192:43:@8101.4]
  wire  _T_23645; // @[LoadQueue.scala 192:43:@8102.4]
  wire  _T_23646; // @[LoadQueue.scala 192:43:@8103.4]
  wire  _T_23647; // @[LoadQueue.scala 192:43:@8104.4]
  wire  _T_23648; // @[LoadQueue.scala 192:43:@8105.4]
  wire  _T_23649; // @[LoadQueue.scala 192:43:@8106.4]
  wire  _T_23650; // @[LoadQueue.scala 192:43:@8107.4]
  wire  _GEN_274; // @[LoadQueue.scala 193:43:@8109.6]
  wire  _GEN_275; // @[LoadQueue.scala 193:43:@8109.6]
  wire  _GEN_276; // @[LoadQueue.scala 193:43:@8109.6]
  wire  _GEN_277; // @[LoadQueue.scala 193:43:@8109.6]
  wire  _GEN_278; // @[LoadQueue.scala 193:43:@8109.6]
  wire  _GEN_279; // @[LoadQueue.scala 193:43:@8109.6]
  wire  _GEN_280; // @[LoadQueue.scala 193:43:@8109.6]
  wire  _GEN_281; // @[LoadQueue.scala 193:43:@8109.6]
  wire  _GEN_283; // @[LoadQueue.scala 194:31:@8110.6]
  wire  _GEN_284; // @[LoadQueue.scala 194:31:@8110.6]
  wire  _GEN_285; // @[LoadQueue.scala 194:31:@8110.6]
  wire  _GEN_286; // @[LoadQueue.scala 194:31:@8110.6]
  wire  _GEN_287; // @[LoadQueue.scala 194:31:@8110.6]
  wire  _GEN_288; // @[LoadQueue.scala 194:31:@8110.6]
  wire  _GEN_289; // @[LoadQueue.scala 194:31:@8110.6]
  wire [31:0] _GEN_291; // @[LoadQueue.scala 195:31:@8111.6]
  wire [31:0] _GEN_292; // @[LoadQueue.scala 195:31:@8111.6]
  wire [31:0] _GEN_293; // @[LoadQueue.scala 195:31:@8111.6]
  wire [31:0] _GEN_294; // @[LoadQueue.scala 195:31:@8111.6]
  wire [31:0] _GEN_295; // @[LoadQueue.scala 195:31:@8111.6]
  wire [31:0] _GEN_296; // @[LoadQueue.scala 195:31:@8111.6]
  wire [31:0] _GEN_297; // @[LoadQueue.scala 195:31:@8111.6]
  wire  lastConflict_1_0; // @[LoadQueue.scala 192:53:@8108.4]
  wire  lastConflict_1_1; // @[LoadQueue.scala 192:53:@8108.4]
  wire  lastConflict_1_2; // @[LoadQueue.scala 192:53:@8108.4]
  wire  lastConflict_1_3; // @[LoadQueue.scala 192:53:@8108.4]
  wire  lastConflict_1_4; // @[LoadQueue.scala 192:53:@8108.4]
  wire  lastConflict_1_5; // @[LoadQueue.scala 192:53:@8108.4]
  wire  lastConflict_1_6; // @[LoadQueue.scala 192:53:@8108.4]
  wire  lastConflict_1_7; // @[LoadQueue.scala 192:53:@8108.4]
  wire  canBypass_1; // @[LoadQueue.scala 192:53:@8108.4]
  wire [31:0] bypassVal_1; // @[LoadQueue.scala 192:53:@8108.4]
  wire [1:0] _T_23716; // @[LoadQueue.scala 191:60:@8141.4]
  wire [1:0] _T_23717; // @[LoadQueue.scala 191:60:@8142.4]
  wire [2:0] _T_23718; // @[LoadQueue.scala 191:60:@8143.4]
  wire [2:0] _T_23719; // @[LoadQueue.scala 191:60:@8144.4]
  wire [2:0] _T_23720; // @[LoadQueue.scala 191:60:@8145.4]
  wire [2:0] _T_23721; // @[LoadQueue.scala 191:60:@8146.4]
  wire  _T_23724; // @[LoadQueue.scala 192:43:@8148.4]
  wire  _T_23725; // @[LoadQueue.scala 192:43:@8149.4]
  wire  _T_23726; // @[LoadQueue.scala 192:43:@8150.4]
  wire  _T_23727; // @[LoadQueue.scala 192:43:@8151.4]
  wire  _T_23728; // @[LoadQueue.scala 192:43:@8152.4]
  wire  _T_23729; // @[LoadQueue.scala 192:43:@8153.4]
  wire  _T_23730; // @[LoadQueue.scala 192:43:@8154.4]
  wire  _GEN_308; // @[LoadQueue.scala 193:43:@8156.6]
  wire  _GEN_309; // @[LoadQueue.scala 193:43:@8156.6]
  wire  _GEN_310; // @[LoadQueue.scala 193:43:@8156.6]
  wire  _GEN_311; // @[LoadQueue.scala 193:43:@8156.6]
  wire  _GEN_312; // @[LoadQueue.scala 193:43:@8156.6]
  wire  _GEN_313; // @[LoadQueue.scala 193:43:@8156.6]
  wire  _GEN_314; // @[LoadQueue.scala 193:43:@8156.6]
  wire  _GEN_315; // @[LoadQueue.scala 193:43:@8156.6]
  wire  _GEN_317; // @[LoadQueue.scala 194:31:@8157.6]
  wire  _GEN_318; // @[LoadQueue.scala 194:31:@8157.6]
  wire  _GEN_319; // @[LoadQueue.scala 194:31:@8157.6]
  wire  _GEN_320; // @[LoadQueue.scala 194:31:@8157.6]
  wire  _GEN_321; // @[LoadQueue.scala 194:31:@8157.6]
  wire  _GEN_322; // @[LoadQueue.scala 194:31:@8157.6]
  wire  _GEN_323; // @[LoadQueue.scala 194:31:@8157.6]
  wire [31:0] _GEN_325; // @[LoadQueue.scala 195:31:@8158.6]
  wire [31:0] _GEN_326; // @[LoadQueue.scala 195:31:@8158.6]
  wire [31:0] _GEN_327; // @[LoadQueue.scala 195:31:@8158.6]
  wire [31:0] _GEN_328; // @[LoadQueue.scala 195:31:@8158.6]
  wire [31:0] _GEN_329; // @[LoadQueue.scala 195:31:@8158.6]
  wire [31:0] _GEN_330; // @[LoadQueue.scala 195:31:@8158.6]
  wire [31:0] _GEN_331; // @[LoadQueue.scala 195:31:@8158.6]
  wire  lastConflict_2_0; // @[LoadQueue.scala 192:53:@8155.4]
  wire  lastConflict_2_1; // @[LoadQueue.scala 192:53:@8155.4]
  wire  lastConflict_2_2; // @[LoadQueue.scala 192:53:@8155.4]
  wire  lastConflict_2_3; // @[LoadQueue.scala 192:53:@8155.4]
  wire  lastConflict_2_4; // @[LoadQueue.scala 192:53:@8155.4]
  wire  lastConflict_2_5; // @[LoadQueue.scala 192:53:@8155.4]
  wire  lastConflict_2_6; // @[LoadQueue.scala 192:53:@8155.4]
  wire  lastConflict_2_7; // @[LoadQueue.scala 192:53:@8155.4]
  wire  canBypass_2; // @[LoadQueue.scala 192:53:@8155.4]
  wire [31:0] bypassVal_2; // @[LoadQueue.scala 192:53:@8155.4]
  wire [1:0] _T_23796; // @[LoadQueue.scala 191:60:@8188.4]
  wire [1:0] _T_23797; // @[LoadQueue.scala 191:60:@8189.4]
  wire [2:0] _T_23798; // @[LoadQueue.scala 191:60:@8190.4]
  wire [2:0] _T_23799; // @[LoadQueue.scala 191:60:@8191.4]
  wire [2:0] _T_23800; // @[LoadQueue.scala 191:60:@8192.4]
  wire [2:0] _T_23801; // @[LoadQueue.scala 191:60:@8193.4]
  wire  _T_23804; // @[LoadQueue.scala 192:43:@8195.4]
  wire  _T_23805; // @[LoadQueue.scala 192:43:@8196.4]
  wire  _T_23806; // @[LoadQueue.scala 192:43:@8197.4]
  wire  _T_23807; // @[LoadQueue.scala 192:43:@8198.4]
  wire  _T_23808; // @[LoadQueue.scala 192:43:@8199.4]
  wire  _T_23809; // @[LoadQueue.scala 192:43:@8200.4]
  wire  _T_23810; // @[LoadQueue.scala 192:43:@8201.4]
  wire  _GEN_342; // @[LoadQueue.scala 193:43:@8203.6]
  wire  _GEN_343; // @[LoadQueue.scala 193:43:@8203.6]
  wire  _GEN_344; // @[LoadQueue.scala 193:43:@8203.6]
  wire  _GEN_345; // @[LoadQueue.scala 193:43:@8203.6]
  wire  _GEN_346; // @[LoadQueue.scala 193:43:@8203.6]
  wire  _GEN_347; // @[LoadQueue.scala 193:43:@8203.6]
  wire  _GEN_348; // @[LoadQueue.scala 193:43:@8203.6]
  wire  _GEN_349; // @[LoadQueue.scala 193:43:@8203.6]
  wire  _GEN_351; // @[LoadQueue.scala 194:31:@8204.6]
  wire  _GEN_352; // @[LoadQueue.scala 194:31:@8204.6]
  wire  _GEN_353; // @[LoadQueue.scala 194:31:@8204.6]
  wire  _GEN_354; // @[LoadQueue.scala 194:31:@8204.6]
  wire  _GEN_355; // @[LoadQueue.scala 194:31:@8204.6]
  wire  _GEN_356; // @[LoadQueue.scala 194:31:@8204.6]
  wire  _GEN_357; // @[LoadQueue.scala 194:31:@8204.6]
  wire [31:0] _GEN_359; // @[LoadQueue.scala 195:31:@8205.6]
  wire [31:0] _GEN_360; // @[LoadQueue.scala 195:31:@8205.6]
  wire [31:0] _GEN_361; // @[LoadQueue.scala 195:31:@8205.6]
  wire [31:0] _GEN_362; // @[LoadQueue.scala 195:31:@8205.6]
  wire [31:0] _GEN_363; // @[LoadQueue.scala 195:31:@8205.6]
  wire [31:0] _GEN_364; // @[LoadQueue.scala 195:31:@8205.6]
  wire [31:0] _GEN_365; // @[LoadQueue.scala 195:31:@8205.6]
  wire  lastConflict_3_0; // @[LoadQueue.scala 192:53:@8202.4]
  wire  lastConflict_3_1; // @[LoadQueue.scala 192:53:@8202.4]
  wire  lastConflict_3_2; // @[LoadQueue.scala 192:53:@8202.4]
  wire  lastConflict_3_3; // @[LoadQueue.scala 192:53:@8202.4]
  wire  lastConflict_3_4; // @[LoadQueue.scala 192:53:@8202.4]
  wire  lastConflict_3_5; // @[LoadQueue.scala 192:53:@8202.4]
  wire  lastConflict_3_6; // @[LoadQueue.scala 192:53:@8202.4]
  wire  lastConflict_3_7; // @[LoadQueue.scala 192:53:@8202.4]
  wire  canBypass_3; // @[LoadQueue.scala 192:53:@8202.4]
  wire [31:0] bypassVal_3; // @[LoadQueue.scala 192:53:@8202.4]
  wire [1:0] _T_23876; // @[LoadQueue.scala 191:60:@8235.4]
  wire [1:0] _T_23877; // @[LoadQueue.scala 191:60:@8236.4]
  wire [2:0] _T_23878; // @[LoadQueue.scala 191:60:@8237.4]
  wire [2:0] _T_23879; // @[LoadQueue.scala 191:60:@8238.4]
  wire [2:0] _T_23880; // @[LoadQueue.scala 191:60:@8239.4]
  wire [2:0] _T_23881; // @[LoadQueue.scala 191:60:@8240.4]
  wire  _T_23884; // @[LoadQueue.scala 192:43:@8242.4]
  wire  _T_23885; // @[LoadQueue.scala 192:43:@8243.4]
  wire  _T_23886; // @[LoadQueue.scala 192:43:@8244.4]
  wire  _T_23887; // @[LoadQueue.scala 192:43:@8245.4]
  wire  _T_23888; // @[LoadQueue.scala 192:43:@8246.4]
  wire  _T_23889; // @[LoadQueue.scala 192:43:@8247.4]
  wire  _T_23890; // @[LoadQueue.scala 192:43:@8248.4]
  wire  _GEN_376; // @[LoadQueue.scala 193:43:@8250.6]
  wire  _GEN_377; // @[LoadQueue.scala 193:43:@8250.6]
  wire  _GEN_378; // @[LoadQueue.scala 193:43:@8250.6]
  wire  _GEN_379; // @[LoadQueue.scala 193:43:@8250.6]
  wire  _GEN_380; // @[LoadQueue.scala 193:43:@8250.6]
  wire  _GEN_381; // @[LoadQueue.scala 193:43:@8250.6]
  wire  _GEN_382; // @[LoadQueue.scala 193:43:@8250.6]
  wire  _GEN_383; // @[LoadQueue.scala 193:43:@8250.6]
  wire  _GEN_385; // @[LoadQueue.scala 194:31:@8251.6]
  wire  _GEN_386; // @[LoadQueue.scala 194:31:@8251.6]
  wire  _GEN_387; // @[LoadQueue.scala 194:31:@8251.6]
  wire  _GEN_388; // @[LoadQueue.scala 194:31:@8251.6]
  wire  _GEN_389; // @[LoadQueue.scala 194:31:@8251.6]
  wire  _GEN_390; // @[LoadQueue.scala 194:31:@8251.6]
  wire  _GEN_391; // @[LoadQueue.scala 194:31:@8251.6]
  wire [31:0] _GEN_393; // @[LoadQueue.scala 195:31:@8252.6]
  wire [31:0] _GEN_394; // @[LoadQueue.scala 195:31:@8252.6]
  wire [31:0] _GEN_395; // @[LoadQueue.scala 195:31:@8252.6]
  wire [31:0] _GEN_396; // @[LoadQueue.scala 195:31:@8252.6]
  wire [31:0] _GEN_397; // @[LoadQueue.scala 195:31:@8252.6]
  wire [31:0] _GEN_398; // @[LoadQueue.scala 195:31:@8252.6]
  wire [31:0] _GEN_399; // @[LoadQueue.scala 195:31:@8252.6]
  wire  lastConflict_4_0; // @[LoadQueue.scala 192:53:@8249.4]
  wire  lastConflict_4_1; // @[LoadQueue.scala 192:53:@8249.4]
  wire  lastConflict_4_2; // @[LoadQueue.scala 192:53:@8249.4]
  wire  lastConflict_4_3; // @[LoadQueue.scala 192:53:@8249.4]
  wire  lastConflict_4_4; // @[LoadQueue.scala 192:53:@8249.4]
  wire  lastConflict_4_5; // @[LoadQueue.scala 192:53:@8249.4]
  wire  lastConflict_4_6; // @[LoadQueue.scala 192:53:@8249.4]
  wire  lastConflict_4_7; // @[LoadQueue.scala 192:53:@8249.4]
  wire  canBypass_4; // @[LoadQueue.scala 192:53:@8249.4]
  wire [31:0] bypassVal_4; // @[LoadQueue.scala 192:53:@8249.4]
  wire [1:0] _T_23956; // @[LoadQueue.scala 191:60:@8282.4]
  wire [1:0] _T_23957; // @[LoadQueue.scala 191:60:@8283.4]
  wire [2:0] _T_23958; // @[LoadQueue.scala 191:60:@8284.4]
  wire [2:0] _T_23959; // @[LoadQueue.scala 191:60:@8285.4]
  wire [2:0] _T_23960; // @[LoadQueue.scala 191:60:@8286.4]
  wire [2:0] _T_23961; // @[LoadQueue.scala 191:60:@8287.4]
  wire  _T_23964; // @[LoadQueue.scala 192:43:@8289.4]
  wire  _T_23965; // @[LoadQueue.scala 192:43:@8290.4]
  wire  _T_23966; // @[LoadQueue.scala 192:43:@8291.4]
  wire  _T_23967; // @[LoadQueue.scala 192:43:@8292.4]
  wire  _T_23968; // @[LoadQueue.scala 192:43:@8293.4]
  wire  _T_23969; // @[LoadQueue.scala 192:43:@8294.4]
  wire  _T_23970; // @[LoadQueue.scala 192:43:@8295.4]
  wire  _GEN_410; // @[LoadQueue.scala 193:43:@8297.6]
  wire  _GEN_411; // @[LoadQueue.scala 193:43:@8297.6]
  wire  _GEN_412; // @[LoadQueue.scala 193:43:@8297.6]
  wire  _GEN_413; // @[LoadQueue.scala 193:43:@8297.6]
  wire  _GEN_414; // @[LoadQueue.scala 193:43:@8297.6]
  wire  _GEN_415; // @[LoadQueue.scala 193:43:@8297.6]
  wire  _GEN_416; // @[LoadQueue.scala 193:43:@8297.6]
  wire  _GEN_417; // @[LoadQueue.scala 193:43:@8297.6]
  wire  _GEN_419; // @[LoadQueue.scala 194:31:@8298.6]
  wire  _GEN_420; // @[LoadQueue.scala 194:31:@8298.6]
  wire  _GEN_421; // @[LoadQueue.scala 194:31:@8298.6]
  wire  _GEN_422; // @[LoadQueue.scala 194:31:@8298.6]
  wire  _GEN_423; // @[LoadQueue.scala 194:31:@8298.6]
  wire  _GEN_424; // @[LoadQueue.scala 194:31:@8298.6]
  wire  _GEN_425; // @[LoadQueue.scala 194:31:@8298.6]
  wire [31:0] _GEN_427; // @[LoadQueue.scala 195:31:@8299.6]
  wire [31:0] _GEN_428; // @[LoadQueue.scala 195:31:@8299.6]
  wire [31:0] _GEN_429; // @[LoadQueue.scala 195:31:@8299.6]
  wire [31:0] _GEN_430; // @[LoadQueue.scala 195:31:@8299.6]
  wire [31:0] _GEN_431; // @[LoadQueue.scala 195:31:@8299.6]
  wire [31:0] _GEN_432; // @[LoadQueue.scala 195:31:@8299.6]
  wire [31:0] _GEN_433; // @[LoadQueue.scala 195:31:@8299.6]
  wire  lastConflict_5_0; // @[LoadQueue.scala 192:53:@8296.4]
  wire  lastConflict_5_1; // @[LoadQueue.scala 192:53:@8296.4]
  wire  lastConflict_5_2; // @[LoadQueue.scala 192:53:@8296.4]
  wire  lastConflict_5_3; // @[LoadQueue.scala 192:53:@8296.4]
  wire  lastConflict_5_4; // @[LoadQueue.scala 192:53:@8296.4]
  wire  lastConflict_5_5; // @[LoadQueue.scala 192:53:@8296.4]
  wire  lastConflict_5_6; // @[LoadQueue.scala 192:53:@8296.4]
  wire  lastConflict_5_7; // @[LoadQueue.scala 192:53:@8296.4]
  wire  canBypass_5; // @[LoadQueue.scala 192:53:@8296.4]
  wire [31:0] bypassVal_5; // @[LoadQueue.scala 192:53:@8296.4]
  wire [1:0] _T_24036; // @[LoadQueue.scala 191:60:@8329.4]
  wire [1:0] _T_24037; // @[LoadQueue.scala 191:60:@8330.4]
  wire [2:0] _T_24038; // @[LoadQueue.scala 191:60:@8331.4]
  wire [2:0] _T_24039; // @[LoadQueue.scala 191:60:@8332.4]
  wire [2:0] _T_24040; // @[LoadQueue.scala 191:60:@8333.4]
  wire [2:0] _T_24041; // @[LoadQueue.scala 191:60:@8334.4]
  wire  _T_24044; // @[LoadQueue.scala 192:43:@8336.4]
  wire  _T_24045; // @[LoadQueue.scala 192:43:@8337.4]
  wire  _T_24046; // @[LoadQueue.scala 192:43:@8338.4]
  wire  _T_24047; // @[LoadQueue.scala 192:43:@8339.4]
  wire  _T_24048; // @[LoadQueue.scala 192:43:@8340.4]
  wire  _T_24049; // @[LoadQueue.scala 192:43:@8341.4]
  wire  _T_24050; // @[LoadQueue.scala 192:43:@8342.4]
  wire  _GEN_444; // @[LoadQueue.scala 193:43:@8344.6]
  wire  _GEN_445; // @[LoadQueue.scala 193:43:@8344.6]
  wire  _GEN_446; // @[LoadQueue.scala 193:43:@8344.6]
  wire  _GEN_447; // @[LoadQueue.scala 193:43:@8344.6]
  wire  _GEN_448; // @[LoadQueue.scala 193:43:@8344.6]
  wire  _GEN_449; // @[LoadQueue.scala 193:43:@8344.6]
  wire  _GEN_450; // @[LoadQueue.scala 193:43:@8344.6]
  wire  _GEN_451; // @[LoadQueue.scala 193:43:@8344.6]
  wire  _GEN_453; // @[LoadQueue.scala 194:31:@8345.6]
  wire  _GEN_454; // @[LoadQueue.scala 194:31:@8345.6]
  wire  _GEN_455; // @[LoadQueue.scala 194:31:@8345.6]
  wire  _GEN_456; // @[LoadQueue.scala 194:31:@8345.6]
  wire  _GEN_457; // @[LoadQueue.scala 194:31:@8345.6]
  wire  _GEN_458; // @[LoadQueue.scala 194:31:@8345.6]
  wire  _GEN_459; // @[LoadQueue.scala 194:31:@8345.6]
  wire [31:0] _GEN_461; // @[LoadQueue.scala 195:31:@8346.6]
  wire [31:0] _GEN_462; // @[LoadQueue.scala 195:31:@8346.6]
  wire [31:0] _GEN_463; // @[LoadQueue.scala 195:31:@8346.6]
  wire [31:0] _GEN_464; // @[LoadQueue.scala 195:31:@8346.6]
  wire [31:0] _GEN_465; // @[LoadQueue.scala 195:31:@8346.6]
  wire [31:0] _GEN_466; // @[LoadQueue.scala 195:31:@8346.6]
  wire [31:0] _GEN_467; // @[LoadQueue.scala 195:31:@8346.6]
  wire  lastConflict_6_0; // @[LoadQueue.scala 192:53:@8343.4]
  wire  lastConflict_6_1; // @[LoadQueue.scala 192:53:@8343.4]
  wire  lastConflict_6_2; // @[LoadQueue.scala 192:53:@8343.4]
  wire  lastConflict_6_3; // @[LoadQueue.scala 192:53:@8343.4]
  wire  lastConflict_6_4; // @[LoadQueue.scala 192:53:@8343.4]
  wire  lastConflict_6_5; // @[LoadQueue.scala 192:53:@8343.4]
  wire  lastConflict_6_6; // @[LoadQueue.scala 192:53:@8343.4]
  wire  lastConflict_6_7; // @[LoadQueue.scala 192:53:@8343.4]
  wire  canBypass_6; // @[LoadQueue.scala 192:53:@8343.4]
  wire [31:0] bypassVal_6; // @[LoadQueue.scala 192:53:@8343.4]
  wire [1:0] _T_24116; // @[LoadQueue.scala 191:60:@8376.4]
  wire [1:0] _T_24117; // @[LoadQueue.scala 191:60:@8377.4]
  wire [2:0] _T_24118; // @[LoadQueue.scala 191:60:@8378.4]
  wire [2:0] _T_24119; // @[LoadQueue.scala 191:60:@8379.4]
  wire [2:0] _T_24120; // @[LoadQueue.scala 191:60:@8380.4]
  wire [2:0] _T_24121; // @[LoadQueue.scala 191:60:@8381.4]
  wire  _T_24124; // @[LoadQueue.scala 192:43:@8383.4]
  wire  _T_24125; // @[LoadQueue.scala 192:43:@8384.4]
  wire  _T_24126; // @[LoadQueue.scala 192:43:@8385.4]
  wire  _T_24127; // @[LoadQueue.scala 192:43:@8386.4]
  wire  _T_24128; // @[LoadQueue.scala 192:43:@8387.4]
  wire  _T_24129; // @[LoadQueue.scala 192:43:@8388.4]
  wire  _T_24130; // @[LoadQueue.scala 192:43:@8389.4]
  wire  _GEN_478; // @[LoadQueue.scala 193:43:@8391.6]
  wire  _GEN_479; // @[LoadQueue.scala 193:43:@8391.6]
  wire  _GEN_480; // @[LoadQueue.scala 193:43:@8391.6]
  wire  _GEN_481; // @[LoadQueue.scala 193:43:@8391.6]
  wire  _GEN_482; // @[LoadQueue.scala 193:43:@8391.6]
  wire  _GEN_483; // @[LoadQueue.scala 193:43:@8391.6]
  wire  _GEN_484; // @[LoadQueue.scala 193:43:@8391.6]
  wire  _GEN_485; // @[LoadQueue.scala 193:43:@8391.6]
  wire  _GEN_487; // @[LoadQueue.scala 194:31:@8392.6]
  wire  _GEN_488; // @[LoadQueue.scala 194:31:@8392.6]
  wire  _GEN_489; // @[LoadQueue.scala 194:31:@8392.6]
  wire  _GEN_490; // @[LoadQueue.scala 194:31:@8392.6]
  wire  _GEN_491; // @[LoadQueue.scala 194:31:@8392.6]
  wire  _GEN_492; // @[LoadQueue.scala 194:31:@8392.6]
  wire  _GEN_493; // @[LoadQueue.scala 194:31:@8392.6]
  wire [31:0] _GEN_495; // @[LoadQueue.scala 195:31:@8393.6]
  wire [31:0] _GEN_496; // @[LoadQueue.scala 195:31:@8393.6]
  wire [31:0] _GEN_497; // @[LoadQueue.scala 195:31:@8393.6]
  wire [31:0] _GEN_498; // @[LoadQueue.scala 195:31:@8393.6]
  wire [31:0] _GEN_499; // @[LoadQueue.scala 195:31:@8393.6]
  wire [31:0] _GEN_500; // @[LoadQueue.scala 195:31:@8393.6]
  wire [31:0] _GEN_501; // @[LoadQueue.scala 195:31:@8393.6]
  wire  lastConflict_7_0; // @[LoadQueue.scala 192:53:@8390.4]
  wire  lastConflict_7_1; // @[LoadQueue.scala 192:53:@8390.4]
  wire  lastConflict_7_2; // @[LoadQueue.scala 192:53:@8390.4]
  wire  lastConflict_7_3; // @[LoadQueue.scala 192:53:@8390.4]
  wire  lastConflict_7_4; // @[LoadQueue.scala 192:53:@8390.4]
  wire  lastConflict_7_5; // @[LoadQueue.scala 192:53:@8390.4]
  wire  lastConflict_7_6; // @[LoadQueue.scala 192:53:@8390.4]
  wire  lastConflict_7_7; // @[LoadQueue.scala 192:53:@8390.4]
  wire  canBypass_7; // @[LoadQueue.scala 192:53:@8390.4]
  wire [31:0] bypassVal_7; // @[LoadQueue.scala 192:53:@8390.4]
  wire [7:0] _T_24174; // @[OneHot.scala 52:12:@8398.4]
  wire  _T_24176; // @[util.scala 33:60:@8400.4]
  wire  _T_24177; // @[util.scala 33:60:@8401.4]
  wire  _T_24178; // @[util.scala 33:60:@8402.4]
  wire  _T_24179; // @[util.scala 33:60:@8403.4]
  wire  _T_24180; // @[util.scala 33:60:@8404.4]
  wire  _T_24181; // @[util.scala 33:60:@8405.4]
  wire  _T_24182; // @[util.scala 33:60:@8406.4]
  wire  _T_24183; // @[util.scala 33:60:@8407.4]
  wire  _T_25168; // @[LoadQueue.scala 229:41:@9154.4]
  wire  _T_25169; // @[LoadQueue.scala 229:38:@9155.4]
  wire  _T_25171; // @[LoadQueue.scala 230:12:@9157.6]
  reg  prevPriorityRequest_7; // @[LoadQueue.scala 207:36:@8716.4]
  reg [31:0] _RAND_243;
  wire  _T_25173; // @[LoadQueue.scala 230:46:@9158.6]
  wire  _T_25174; // @[LoadQueue.scala 230:43:@9159.6]
  wire  _T_25176; // @[LoadQueue.scala 230:84:@9160.6]
  wire  _T_25177; // @[LoadQueue.scala 230:81:@9161.6]
  wire  _T_25180; // @[LoadQueue.scala 233:86:@9164.8]
  wire  _T_25181; // @[LoadQueue.scala 233:86:@9165.8]
  wire  _T_25182; // @[LoadQueue.scala 233:86:@9166.8]
  wire  _T_25183; // @[LoadQueue.scala 233:86:@9167.8]
  wire  _T_25184; // @[LoadQueue.scala 233:86:@9168.8]
  wire  _T_25185; // @[LoadQueue.scala 233:86:@9169.8]
  wire  _T_25186; // @[LoadQueue.scala 233:86:@9170.8]
  wire  _T_25188; // @[LoadQueue.scala 233:38:@9171.8]
  wire  _T_25199; // @[LoadQueue.scala 234:11:@9180.8]
  wire  _T_25200; // @[LoadQueue.scala 233:103:@9181.8]
  wire  _GEN_564; // @[LoadQueue.scala 230:110:@9162.6]
  wire  loadRequest_7; // @[LoadQueue.scala 229:71:@9156.4]
  wire [7:0] _T_24208; // @[Mux.scala 31:69:@8417.4]
  wire  _T_25116; // @[LoadQueue.scala 229:41:@9104.4]
  wire  _T_25117; // @[LoadQueue.scala 229:38:@9105.4]
  wire  _T_25119; // @[LoadQueue.scala 230:12:@9107.6]
  reg  prevPriorityRequest_6; // @[LoadQueue.scala 207:36:@8716.4]
  reg [31:0] _RAND_244;
  wire  _T_25121; // @[LoadQueue.scala 230:46:@9108.6]
  wire  _T_25122; // @[LoadQueue.scala 230:43:@9109.6]
  wire  _T_25124; // @[LoadQueue.scala 230:84:@9110.6]
  wire  _T_25125; // @[LoadQueue.scala 230:81:@9111.6]
  wire  _T_25128; // @[LoadQueue.scala 233:86:@9114.8]
  wire  _T_25129; // @[LoadQueue.scala 233:86:@9115.8]
  wire  _T_25130; // @[LoadQueue.scala 233:86:@9116.8]
  wire  _T_25131; // @[LoadQueue.scala 233:86:@9117.8]
  wire  _T_25132; // @[LoadQueue.scala 233:86:@9118.8]
  wire  _T_25133; // @[LoadQueue.scala 233:86:@9119.8]
  wire  _T_25134; // @[LoadQueue.scala 233:86:@9120.8]
  wire  _T_25136; // @[LoadQueue.scala 233:38:@9121.8]
  wire  _T_25147; // @[LoadQueue.scala 234:11:@9130.8]
  wire  _T_25148; // @[LoadQueue.scala 233:103:@9131.8]
  wire  _GEN_560; // @[LoadQueue.scala 230:110:@9112.6]
  wire  loadRequest_6; // @[LoadQueue.scala 229:71:@9106.4]
  wire [7:0] _T_24209; // @[Mux.scala 31:69:@8418.4]
  wire  _T_25064; // @[LoadQueue.scala 229:41:@9054.4]
  wire  _T_25065; // @[LoadQueue.scala 229:38:@9055.4]
  wire  _T_25067; // @[LoadQueue.scala 230:12:@9057.6]
  reg  prevPriorityRequest_5; // @[LoadQueue.scala 207:36:@8716.4]
  reg [31:0] _RAND_245;
  wire  _T_25069; // @[LoadQueue.scala 230:46:@9058.6]
  wire  _T_25070; // @[LoadQueue.scala 230:43:@9059.6]
  wire  _T_25072; // @[LoadQueue.scala 230:84:@9060.6]
  wire  _T_25073; // @[LoadQueue.scala 230:81:@9061.6]
  wire  _T_25076; // @[LoadQueue.scala 233:86:@9064.8]
  wire  _T_25077; // @[LoadQueue.scala 233:86:@9065.8]
  wire  _T_25078; // @[LoadQueue.scala 233:86:@9066.8]
  wire  _T_25079; // @[LoadQueue.scala 233:86:@9067.8]
  wire  _T_25080; // @[LoadQueue.scala 233:86:@9068.8]
  wire  _T_25081; // @[LoadQueue.scala 233:86:@9069.8]
  wire  _T_25082; // @[LoadQueue.scala 233:86:@9070.8]
  wire  _T_25084; // @[LoadQueue.scala 233:38:@9071.8]
  wire  _T_25095; // @[LoadQueue.scala 234:11:@9080.8]
  wire  _T_25096; // @[LoadQueue.scala 233:103:@9081.8]
  wire  _GEN_556; // @[LoadQueue.scala 230:110:@9062.6]
  wire  loadRequest_5; // @[LoadQueue.scala 229:71:@9056.4]
  wire [7:0] _T_24210; // @[Mux.scala 31:69:@8419.4]
  wire  _T_25012; // @[LoadQueue.scala 229:41:@9004.4]
  wire  _T_25013; // @[LoadQueue.scala 229:38:@9005.4]
  wire  _T_25015; // @[LoadQueue.scala 230:12:@9007.6]
  reg  prevPriorityRequest_4; // @[LoadQueue.scala 207:36:@8716.4]
  reg [31:0] _RAND_246;
  wire  _T_25017; // @[LoadQueue.scala 230:46:@9008.6]
  wire  _T_25018; // @[LoadQueue.scala 230:43:@9009.6]
  wire  _T_25020; // @[LoadQueue.scala 230:84:@9010.6]
  wire  _T_25021; // @[LoadQueue.scala 230:81:@9011.6]
  wire  _T_25024; // @[LoadQueue.scala 233:86:@9014.8]
  wire  _T_25025; // @[LoadQueue.scala 233:86:@9015.8]
  wire  _T_25026; // @[LoadQueue.scala 233:86:@9016.8]
  wire  _T_25027; // @[LoadQueue.scala 233:86:@9017.8]
  wire  _T_25028; // @[LoadQueue.scala 233:86:@9018.8]
  wire  _T_25029; // @[LoadQueue.scala 233:86:@9019.8]
  wire  _T_25030; // @[LoadQueue.scala 233:86:@9020.8]
  wire  _T_25032; // @[LoadQueue.scala 233:38:@9021.8]
  wire  _T_25043; // @[LoadQueue.scala 234:11:@9030.8]
  wire  _T_25044; // @[LoadQueue.scala 233:103:@9031.8]
  wire  _GEN_552; // @[LoadQueue.scala 230:110:@9012.6]
  wire  loadRequest_4; // @[LoadQueue.scala 229:71:@9006.4]
  wire [7:0] _T_24211; // @[Mux.scala 31:69:@8420.4]
  wire  _T_24960; // @[LoadQueue.scala 229:41:@8954.4]
  wire  _T_24961; // @[LoadQueue.scala 229:38:@8955.4]
  wire  _T_24963; // @[LoadQueue.scala 230:12:@8957.6]
  reg  prevPriorityRequest_3; // @[LoadQueue.scala 207:36:@8716.4]
  reg [31:0] _RAND_247;
  wire  _T_24965; // @[LoadQueue.scala 230:46:@8958.6]
  wire  _T_24966; // @[LoadQueue.scala 230:43:@8959.6]
  wire  _T_24968; // @[LoadQueue.scala 230:84:@8960.6]
  wire  _T_24969; // @[LoadQueue.scala 230:81:@8961.6]
  wire  _T_24972; // @[LoadQueue.scala 233:86:@8964.8]
  wire  _T_24973; // @[LoadQueue.scala 233:86:@8965.8]
  wire  _T_24974; // @[LoadQueue.scala 233:86:@8966.8]
  wire  _T_24975; // @[LoadQueue.scala 233:86:@8967.8]
  wire  _T_24976; // @[LoadQueue.scala 233:86:@8968.8]
  wire  _T_24977; // @[LoadQueue.scala 233:86:@8969.8]
  wire  _T_24978; // @[LoadQueue.scala 233:86:@8970.8]
  wire  _T_24980; // @[LoadQueue.scala 233:38:@8971.8]
  wire  _T_24991; // @[LoadQueue.scala 234:11:@8980.8]
  wire  _T_24992; // @[LoadQueue.scala 233:103:@8981.8]
  wire  _GEN_548; // @[LoadQueue.scala 230:110:@8962.6]
  wire  loadRequest_3; // @[LoadQueue.scala 229:71:@8956.4]
  wire [7:0] _T_24212; // @[Mux.scala 31:69:@8421.4]
  wire  _T_24908; // @[LoadQueue.scala 229:41:@8904.4]
  wire  _T_24909; // @[LoadQueue.scala 229:38:@8905.4]
  wire  _T_24911; // @[LoadQueue.scala 230:12:@8907.6]
  reg  prevPriorityRequest_2; // @[LoadQueue.scala 207:36:@8716.4]
  reg [31:0] _RAND_248;
  wire  _T_24913; // @[LoadQueue.scala 230:46:@8908.6]
  wire  _T_24914; // @[LoadQueue.scala 230:43:@8909.6]
  wire  _T_24916; // @[LoadQueue.scala 230:84:@8910.6]
  wire  _T_24917; // @[LoadQueue.scala 230:81:@8911.6]
  wire  _T_24920; // @[LoadQueue.scala 233:86:@8914.8]
  wire  _T_24921; // @[LoadQueue.scala 233:86:@8915.8]
  wire  _T_24922; // @[LoadQueue.scala 233:86:@8916.8]
  wire  _T_24923; // @[LoadQueue.scala 233:86:@8917.8]
  wire  _T_24924; // @[LoadQueue.scala 233:86:@8918.8]
  wire  _T_24925; // @[LoadQueue.scala 233:86:@8919.8]
  wire  _T_24926; // @[LoadQueue.scala 233:86:@8920.8]
  wire  _T_24928; // @[LoadQueue.scala 233:38:@8921.8]
  wire  _T_24939; // @[LoadQueue.scala 234:11:@8930.8]
  wire  _T_24940; // @[LoadQueue.scala 233:103:@8931.8]
  wire  _GEN_544; // @[LoadQueue.scala 230:110:@8912.6]
  wire  loadRequest_2; // @[LoadQueue.scala 229:71:@8906.4]
  wire [7:0] _T_24213; // @[Mux.scala 31:69:@8422.4]
  wire  _T_24856; // @[LoadQueue.scala 229:41:@8854.4]
  wire  _T_24857; // @[LoadQueue.scala 229:38:@8855.4]
  wire  _T_24859; // @[LoadQueue.scala 230:12:@8857.6]
  reg  prevPriorityRequest_1; // @[LoadQueue.scala 207:36:@8716.4]
  reg [31:0] _RAND_249;
  wire  _T_24861; // @[LoadQueue.scala 230:46:@8858.6]
  wire  _T_24862; // @[LoadQueue.scala 230:43:@8859.6]
  wire  _T_24864; // @[LoadQueue.scala 230:84:@8860.6]
  wire  _T_24865; // @[LoadQueue.scala 230:81:@8861.6]
  wire  _T_24868; // @[LoadQueue.scala 233:86:@8864.8]
  wire  _T_24869; // @[LoadQueue.scala 233:86:@8865.8]
  wire  _T_24870; // @[LoadQueue.scala 233:86:@8866.8]
  wire  _T_24871; // @[LoadQueue.scala 233:86:@8867.8]
  wire  _T_24872; // @[LoadQueue.scala 233:86:@8868.8]
  wire  _T_24873; // @[LoadQueue.scala 233:86:@8869.8]
  wire  _T_24874; // @[LoadQueue.scala 233:86:@8870.8]
  wire  _T_24876; // @[LoadQueue.scala 233:38:@8871.8]
  wire  _T_24887; // @[LoadQueue.scala 234:11:@8880.8]
  wire  _T_24888; // @[LoadQueue.scala 233:103:@8881.8]
  wire  _GEN_540; // @[LoadQueue.scala 230:110:@8862.6]
  wire  loadRequest_1; // @[LoadQueue.scala 229:71:@8856.4]
  wire [7:0] _T_24214; // @[Mux.scala 31:69:@8423.4]
  wire  _T_24804; // @[LoadQueue.scala 229:41:@8804.4]
  wire  _T_24805; // @[LoadQueue.scala 229:38:@8805.4]
  wire  _T_24807; // @[LoadQueue.scala 230:12:@8807.6]
  reg  prevPriorityRequest_0; // @[LoadQueue.scala 207:36:@8716.4]
  reg [31:0] _RAND_250;
  wire  _T_24809; // @[LoadQueue.scala 230:46:@8808.6]
  wire  _T_24810; // @[LoadQueue.scala 230:43:@8809.6]
  wire  _T_24812; // @[LoadQueue.scala 230:84:@8810.6]
  wire  _T_24813; // @[LoadQueue.scala 230:81:@8811.6]
  wire  _T_24816; // @[LoadQueue.scala 233:86:@8814.8]
  wire  _T_24817; // @[LoadQueue.scala 233:86:@8815.8]
  wire  _T_24818; // @[LoadQueue.scala 233:86:@8816.8]
  wire  _T_24819; // @[LoadQueue.scala 233:86:@8817.8]
  wire  _T_24820; // @[LoadQueue.scala 233:86:@8818.8]
  wire  _T_24821; // @[LoadQueue.scala 233:86:@8819.8]
  wire  _T_24822; // @[LoadQueue.scala 233:86:@8820.8]
  wire  _T_24824; // @[LoadQueue.scala 233:38:@8821.8]
  wire  _T_24835; // @[LoadQueue.scala 234:11:@8830.8]
  wire  _T_24836; // @[LoadQueue.scala 233:103:@8831.8]
  wire  _GEN_536; // @[LoadQueue.scala 230:110:@8812.6]
  wire  loadRequest_0; // @[LoadQueue.scala 229:71:@8806.4]
  wire [7:0] _T_24215; // @[Mux.scala 31:69:@8424.4]
  wire  _T_24216; // @[OneHot.scala 66:30:@8425.4]
  wire  _T_24217; // @[OneHot.scala 66:30:@8426.4]
  wire  _T_24218; // @[OneHot.scala 66:30:@8427.4]
  wire  _T_24219; // @[OneHot.scala 66:30:@8428.4]
  wire  _T_24220; // @[OneHot.scala 66:30:@8429.4]
  wire  _T_24221; // @[OneHot.scala 66:30:@8430.4]
  wire  _T_24222; // @[OneHot.scala 66:30:@8431.4]
  wire  _T_24223; // @[OneHot.scala 66:30:@8432.4]
  wire [7:0] _T_24248; // @[Mux.scala 31:69:@8442.4]
  wire [7:0] _T_24249; // @[Mux.scala 31:69:@8443.4]
  wire [7:0] _T_24250; // @[Mux.scala 31:69:@8444.4]
  wire [7:0] _T_24251; // @[Mux.scala 31:69:@8445.4]
  wire [7:0] _T_24252; // @[Mux.scala 31:69:@8446.4]
  wire [7:0] _T_24253; // @[Mux.scala 31:69:@8447.4]
  wire [7:0] _T_24254; // @[Mux.scala 31:69:@8448.4]
  wire [7:0] _T_24255; // @[Mux.scala 31:69:@8449.4]
  wire  _T_24256; // @[OneHot.scala 66:30:@8450.4]
  wire  _T_24257; // @[OneHot.scala 66:30:@8451.4]
  wire  _T_24258; // @[OneHot.scala 66:30:@8452.4]
  wire  _T_24259; // @[OneHot.scala 66:30:@8453.4]
  wire  _T_24260; // @[OneHot.scala 66:30:@8454.4]
  wire  _T_24261; // @[OneHot.scala 66:30:@8455.4]
  wire  _T_24262; // @[OneHot.scala 66:30:@8456.4]
  wire  _T_24263; // @[OneHot.scala 66:30:@8457.4]
  wire [7:0] _T_24288; // @[Mux.scala 31:69:@8467.4]
  wire [7:0] _T_24289; // @[Mux.scala 31:69:@8468.4]
  wire [7:0] _T_24290; // @[Mux.scala 31:69:@8469.4]
  wire [7:0] _T_24291; // @[Mux.scala 31:69:@8470.4]
  wire [7:0] _T_24292; // @[Mux.scala 31:69:@8471.4]
  wire [7:0] _T_24293; // @[Mux.scala 31:69:@8472.4]
  wire [7:0] _T_24294; // @[Mux.scala 31:69:@8473.4]
  wire [7:0] _T_24295; // @[Mux.scala 31:69:@8474.4]
  wire  _T_24296; // @[OneHot.scala 66:30:@8475.4]
  wire  _T_24297; // @[OneHot.scala 66:30:@8476.4]
  wire  _T_24298; // @[OneHot.scala 66:30:@8477.4]
  wire  _T_24299; // @[OneHot.scala 66:30:@8478.4]
  wire  _T_24300; // @[OneHot.scala 66:30:@8479.4]
  wire  _T_24301; // @[OneHot.scala 66:30:@8480.4]
  wire  _T_24302; // @[OneHot.scala 66:30:@8481.4]
  wire  _T_24303; // @[OneHot.scala 66:30:@8482.4]
  wire [7:0] _T_24328; // @[Mux.scala 31:69:@8492.4]
  wire [7:0] _T_24329; // @[Mux.scala 31:69:@8493.4]
  wire [7:0] _T_24330; // @[Mux.scala 31:69:@8494.4]
  wire [7:0] _T_24331; // @[Mux.scala 31:69:@8495.4]
  wire [7:0] _T_24332; // @[Mux.scala 31:69:@8496.4]
  wire [7:0] _T_24333; // @[Mux.scala 31:69:@8497.4]
  wire [7:0] _T_24334; // @[Mux.scala 31:69:@8498.4]
  wire [7:0] _T_24335; // @[Mux.scala 31:69:@8499.4]
  wire  _T_24336; // @[OneHot.scala 66:30:@8500.4]
  wire  _T_24337; // @[OneHot.scala 66:30:@8501.4]
  wire  _T_24338; // @[OneHot.scala 66:30:@8502.4]
  wire  _T_24339; // @[OneHot.scala 66:30:@8503.4]
  wire  _T_24340; // @[OneHot.scala 66:30:@8504.4]
  wire  _T_24341; // @[OneHot.scala 66:30:@8505.4]
  wire  _T_24342; // @[OneHot.scala 66:30:@8506.4]
  wire  _T_24343; // @[OneHot.scala 66:30:@8507.4]
  wire [7:0] _T_24368; // @[Mux.scala 31:69:@8517.4]
  wire [7:0] _T_24369; // @[Mux.scala 31:69:@8518.4]
  wire [7:0] _T_24370; // @[Mux.scala 31:69:@8519.4]
  wire [7:0] _T_24371; // @[Mux.scala 31:69:@8520.4]
  wire [7:0] _T_24372; // @[Mux.scala 31:69:@8521.4]
  wire [7:0] _T_24373; // @[Mux.scala 31:69:@8522.4]
  wire [7:0] _T_24374; // @[Mux.scala 31:69:@8523.4]
  wire [7:0] _T_24375; // @[Mux.scala 31:69:@8524.4]
  wire  _T_24376; // @[OneHot.scala 66:30:@8525.4]
  wire  _T_24377; // @[OneHot.scala 66:30:@8526.4]
  wire  _T_24378; // @[OneHot.scala 66:30:@8527.4]
  wire  _T_24379; // @[OneHot.scala 66:30:@8528.4]
  wire  _T_24380; // @[OneHot.scala 66:30:@8529.4]
  wire  _T_24381; // @[OneHot.scala 66:30:@8530.4]
  wire  _T_24382; // @[OneHot.scala 66:30:@8531.4]
  wire  _T_24383; // @[OneHot.scala 66:30:@8532.4]
  wire [7:0] _T_24408; // @[Mux.scala 31:69:@8542.4]
  wire [7:0] _T_24409; // @[Mux.scala 31:69:@8543.4]
  wire [7:0] _T_24410; // @[Mux.scala 31:69:@8544.4]
  wire [7:0] _T_24411; // @[Mux.scala 31:69:@8545.4]
  wire [7:0] _T_24412; // @[Mux.scala 31:69:@8546.4]
  wire [7:0] _T_24413; // @[Mux.scala 31:69:@8547.4]
  wire [7:0] _T_24414; // @[Mux.scala 31:69:@8548.4]
  wire [7:0] _T_24415; // @[Mux.scala 31:69:@8549.4]
  wire  _T_24416; // @[OneHot.scala 66:30:@8550.4]
  wire  _T_24417; // @[OneHot.scala 66:30:@8551.4]
  wire  _T_24418; // @[OneHot.scala 66:30:@8552.4]
  wire  _T_24419; // @[OneHot.scala 66:30:@8553.4]
  wire  _T_24420; // @[OneHot.scala 66:30:@8554.4]
  wire  _T_24421; // @[OneHot.scala 66:30:@8555.4]
  wire  _T_24422; // @[OneHot.scala 66:30:@8556.4]
  wire  _T_24423; // @[OneHot.scala 66:30:@8557.4]
  wire [7:0] _T_24448; // @[Mux.scala 31:69:@8567.4]
  wire [7:0] _T_24449; // @[Mux.scala 31:69:@8568.4]
  wire [7:0] _T_24450; // @[Mux.scala 31:69:@8569.4]
  wire [7:0] _T_24451; // @[Mux.scala 31:69:@8570.4]
  wire [7:0] _T_24452; // @[Mux.scala 31:69:@8571.4]
  wire [7:0] _T_24453; // @[Mux.scala 31:69:@8572.4]
  wire [7:0] _T_24454; // @[Mux.scala 31:69:@8573.4]
  wire [7:0] _T_24455; // @[Mux.scala 31:69:@8574.4]
  wire  _T_24456; // @[OneHot.scala 66:30:@8575.4]
  wire  _T_24457; // @[OneHot.scala 66:30:@8576.4]
  wire  _T_24458; // @[OneHot.scala 66:30:@8577.4]
  wire  _T_24459; // @[OneHot.scala 66:30:@8578.4]
  wire  _T_24460; // @[OneHot.scala 66:30:@8579.4]
  wire  _T_24461; // @[OneHot.scala 66:30:@8580.4]
  wire  _T_24462; // @[OneHot.scala 66:30:@8581.4]
  wire  _T_24463; // @[OneHot.scala 66:30:@8582.4]
  wire [7:0] _T_24488; // @[Mux.scala 31:69:@8592.4]
  wire [7:0] _T_24489; // @[Mux.scala 31:69:@8593.4]
  wire [7:0] _T_24490; // @[Mux.scala 31:69:@8594.4]
  wire [7:0] _T_24491; // @[Mux.scala 31:69:@8595.4]
  wire [7:0] _T_24492; // @[Mux.scala 31:69:@8596.4]
  wire [7:0] _T_24493; // @[Mux.scala 31:69:@8597.4]
  wire [7:0] _T_24494; // @[Mux.scala 31:69:@8598.4]
  wire [7:0] _T_24495; // @[Mux.scala 31:69:@8599.4]
  wire  _T_24496; // @[OneHot.scala 66:30:@8600.4]
  wire  _T_24497; // @[OneHot.scala 66:30:@8601.4]
  wire  _T_24498; // @[OneHot.scala 66:30:@8602.4]
  wire  _T_24499; // @[OneHot.scala 66:30:@8603.4]
  wire  _T_24500; // @[OneHot.scala 66:30:@8604.4]
  wire  _T_24501; // @[OneHot.scala 66:30:@8605.4]
  wire  _T_24502; // @[OneHot.scala 66:30:@8606.4]
  wire  _T_24503; // @[OneHot.scala 66:30:@8607.4]
  wire [7:0] _T_24544; // @[Mux.scala 19:72:@8623.4]
  wire [7:0] _T_24546; // @[Mux.scala 19:72:@8624.4]
  wire [7:0] _T_24553; // @[Mux.scala 19:72:@8631.4]
  wire [7:0] _T_24555; // @[Mux.scala 19:72:@8632.4]
  wire [7:0] _T_24562; // @[Mux.scala 19:72:@8639.4]
  wire [7:0] _T_24564; // @[Mux.scala 19:72:@8640.4]
  wire [7:0] _T_24571; // @[Mux.scala 19:72:@8647.4]
  wire [7:0] _T_24573; // @[Mux.scala 19:72:@8648.4]
  wire [7:0] _T_24580; // @[Mux.scala 19:72:@8655.4]
  wire [7:0] _T_24582; // @[Mux.scala 19:72:@8656.4]
  wire [7:0] _T_24589; // @[Mux.scala 19:72:@8663.4]
  wire [7:0] _T_24591; // @[Mux.scala 19:72:@8664.4]
  wire [7:0] _T_24598; // @[Mux.scala 19:72:@8671.4]
  wire [7:0] _T_24600; // @[Mux.scala 19:72:@8672.4]
  wire [7:0] _T_24607; // @[Mux.scala 19:72:@8679.4]
  wire [7:0] _T_24609; // @[Mux.scala 19:72:@8680.4]
  wire [7:0] _T_24610; // @[Mux.scala 19:72:@8681.4]
  wire [7:0] _T_24611; // @[Mux.scala 19:72:@8682.4]
  wire [7:0] _T_24612; // @[Mux.scala 19:72:@8683.4]
  wire [7:0] _T_24613; // @[Mux.scala 19:72:@8684.4]
  wire [7:0] _T_24614; // @[Mux.scala 19:72:@8685.4]
  wire [7:0] _T_24615; // @[Mux.scala 19:72:@8686.4]
  wire [7:0] _T_24616; // @[Mux.scala 19:72:@8687.4]
  wire  priorityLoadRequest_0; // @[Mux.scala 19:72:@8691.4]
  wire  priorityLoadRequest_1; // @[Mux.scala 19:72:@8693.4]
  wire  priorityLoadRequest_2; // @[Mux.scala 19:72:@8695.4]
  wire  priorityLoadRequest_3; // @[Mux.scala 19:72:@8697.4]
  wire  priorityLoadRequest_4; // @[Mux.scala 19:72:@8699.4]
  wire  priorityLoadRequest_5; // @[Mux.scala 19:72:@8701.4]
  wire  priorityLoadRequest_6; // @[Mux.scala 19:72:@8703.4]
  wire  priorityLoadRequest_7; // @[Mux.scala 19:72:@8705.4]
  wire  _GEN_512; // @[LoadQueue.scala 208:31:@8717.4]
  wire  _GEN_513; // @[LoadQueue.scala 208:31:@8717.4]
  wire  _GEN_514; // @[LoadQueue.scala 208:31:@8717.4]
  wire  _GEN_515; // @[LoadQueue.scala 208:31:@8717.4]
  wire  _GEN_516; // @[LoadQueue.scala 208:31:@8717.4]
  wire  _GEN_517; // @[LoadQueue.scala 208:31:@8717.4]
  wire  _GEN_518; // @[LoadQueue.scala 208:31:@8717.4]
  wire  _GEN_519; // @[LoadQueue.scala 208:31:@8717.4]
  wire [7:0] _T_24843; // @[LoadQueue.scala 238:58:@8839.8]
  wire [7:0] _T_24850; // @[LoadQueue.scala 238:96:@8846.8]
  wire  _T_24851; // @[LoadQueue.scala 238:61:@8847.8]
  wire  _T_24852; // @[LoadQueue.scala 237:64:@8848.8]
  wire  _GEN_537; // @[LoadQueue.scala 230:110:@8812.6]
  wire  bypassRequest_0; // @[LoadQueue.scala 229:71:@8806.4]
  wire  _GEN_520; // @[LoadQueue.scala 217:34:@8750.6]
  wire  _GEN_521; // @[LoadQueue.scala 215:23:@8746.4]
  wire [7:0] _T_24895; // @[LoadQueue.scala 238:58:@8889.8]
  wire [7:0] _T_24902; // @[LoadQueue.scala 238:96:@8896.8]
  wire  _T_24903; // @[LoadQueue.scala 238:61:@8897.8]
  wire  _T_24904; // @[LoadQueue.scala 237:64:@8898.8]
  wire  _GEN_541; // @[LoadQueue.scala 230:110:@8862.6]
  wire  bypassRequest_1; // @[LoadQueue.scala 229:71:@8856.4]
  wire  _GEN_522; // @[LoadQueue.scala 217:34:@8757.6]
  wire  _GEN_523; // @[LoadQueue.scala 215:23:@8753.4]
  wire [7:0] _T_24947; // @[LoadQueue.scala 238:58:@8939.8]
  wire [7:0] _T_24954; // @[LoadQueue.scala 238:96:@8946.8]
  wire  _T_24955; // @[LoadQueue.scala 238:61:@8947.8]
  wire  _T_24956; // @[LoadQueue.scala 237:64:@8948.8]
  wire  _GEN_545; // @[LoadQueue.scala 230:110:@8912.6]
  wire  bypassRequest_2; // @[LoadQueue.scala 229:71:@8906.4]
  wire  _GEN_524; // @[LoadQueue.scala 217:34:@8764.6]
  wire  _GEN_525; // @[LoadQueue.scala 215:23:@8760.4]
  wire [7:0] _T_24999; // @[LoadQueue.scala 238:58:@8989.8]
  wire [7:0] _T_25006; // @[LoadQueue.scala 238:96:@8996.8]
  wire  _T_25007; // @[LoadQueue.scala 238:61:@8997.8]
  wire  _T_25008; // @[LoadQueue.scala 237:64:@8998.8]
  wire  _GEN_549; // @[LoadQueue.scala 230:110:@8962.6]
  wire  bypassRequest_3; // @[LoadQueue.scala 229:71:@8956.4]
  wire  _GEN_526; // @[LoadQueue.scala 217:34:@8771.6]
  wire  _GEN_527; // @[LoadQueue.scala 215:23:@8767.4]
  wire [7:0] _T_25051; // @[LoadQueue.scala 238:58:@9039.8]
  wire [7:0] _T_25058; // @[LoadQueue.scala 238:96:@9046.8]
  wire  _T_25059; // @[LoadQueue.scala 238:61:@9047.8]
  wire  _T_25060; // @[LoadQueue.scala 237:64:@9048.8]
  wire  _GEN_553; // @[LoadQueue.scala 230:110:@9012.6]
  wire  bypassRequest_4; // @[LoadQueue.scala 229:71:@9006.4]
  wire  _GEN_528; // @[LoadQueue.scala 217:34:@8778.6]
  wire  _GEN_529; // @[LoadQueue.scala 215:23:@8774.4]
  wire [7:0] _T_25103; // @[LoadQueue.scala 238:58:@9089.8]
  wire [7:0] _T_25110; // @[LoadQueue.scala 238:96:@9096.8]
  wire  _T_25111; // @[LoadQueue.scala 238:61:@9097.8]
  wire  _T_25112; // @[LoadQueue.scala 237:64:@9098.8]
  wire  _GEN_557; // @[LoadQueue.scala 230:110:@9062.6]
  wire  bypassRequest_5; // @[LoadQueue.scala 229:71:@9056.4]
  wire  _GEN_530; // @[LoadQueue.scala 217:34:@8785.6]
  wire  _GEN_531; // @[LoadQueue.scala 215:23:@8781.4]
  wire [7:0] _T_25155; // @[LoadQueue.scala 238:58:@9139.8]
  wire [7:0] _T_25162; // @[LoadQueue.scala 238:96:@9146.8]
  wire  _T_25163; // @[LoadQueue.scala 238:61:@9147.8]
  wire  _T_25164; // @[LoadQueue.scala 237:64:@9148.8]
  wire  _GEN_561; // @[LoadQueue.scala 230:110:@9112.6]
  wire  bypassRequest_6; // @[LoadQueue.scala 229:71:@9106.4]
  wire  _GEN_532; // @[LoadQueue.scala 217:34:@8792.6]
  wire  _GEN_533; // @[LoadQueue.scala 215:23:@8788.4]
  wire [7:0] _T_25207; // @[LoadQueue.scala 238:58:@9189.8]
  wire [7:0] _T_25214; // @[LoadQueue.scala 238:96:@9196.8]
  wire  _T_25215; // @[LoadQueue.scala 238:61:@9197.8]
  wire  _T_25216; // @[LoadQueue.scala 237:64:@9198.8]
  wire  _GEN_565; // @[LoadQueue.scala 230:110:@9162.6]
  wire  bypassRequest_7; // @[LoadQueue.scala 229:71:@9156.4]
  wire  _GEN_534; // @[LoadQueue.scala 217:34:@8799.6]
  wire  _GEN_535; // @[LoadQueue.scala 215:23:@8795.4]
  wire  _T_25220; // @[LoadQueue.scala 247:28:@9204.4]
  wire  _T_25221; // @[LoadQueue.scala 247:28:@9205.4]
  wire  _T_25222; // @[LoadQueue.scala 247:28:@9206.4]
  wire  _T_25223; // @[LoadQueue.scala 247:28:@9207.4]
  wire  _T_25224; // @[LoadQueue.scala 247:28:@9208.4]
  wire  _T_25225; // @[LoadQueue.scala 247:28:@9209.4]
  wire  _T_25226; // @[LoadQueue.scala 247:28:@9210.4]
  wire [2:0] _T_25235; // @[Mux.scala 31:69:@9212.6]
  wire [2:0] _T_25236; // @[Mux.scala 31:69:@9213.6]
  wire [2:0] _T_25237; // @[Mux.scala 31:69:@9214.6]
  wire [2:0] _T_25238; // @[Mux.scala 31:69:@9215.6]
  wire [2:0] _T_25239; // @[Mux.scala 31:69:@9216.6]
  wire [2:0] _T_25240; // @[Mux.scala 31:69:@9217.6]
  wire [2:0] _T_25241; // @[Mux.scala 31:69:@9218.6]
  wire [31:0] _GEN_569; // @[LoadQueue.scala 248:24:@9219.6]
  wire [31:0] _GEN_570; // @[LoadQueue.scala 248:24:@9219.6]
  wire [31:0] _GEN_571; // @[LoadQueue.scala 248:24:@9219.6]
  wire [31:0] _GEN_572; // @[LoadQueue.scala 248:24:@9219.6]
  wire [31:0] _GEN_573; // @[LoadQueue.scala 248:24:@9219.6]
  wire [31:0] _GEN_574; // @[LoadQueue.scala 248:24:@9219.6]
  wire [31:0] _GEN_575; // @[LoadQueue.scala 248:24:@9219.6]
  wire  _T_25249; // @[LoadQueue.scala 261:41:@9230.6]
  wire  _GEN_578; // @[LoadQueue.scala 261:62:@9231.6]
  wire  _GEN_579; // @[LoadQueue.scala 259:25:@9226.4]
  wire  _T_25252; // @[LoadQueue.scala 261:41:@9238.6]
  wire  _GEN_580; // @[LoadQueue.scala 261:62:@9239.6]
  wire  _GEN_581; // @[LoadQueue.scala 259:25:@9234.4]
  wire  _T_25255; // @[LoadQueue.scala 261:41:@9246.6]
  wire  _GEN_582; // @[LoadQueue.scala 261:62:@9247.6]
  wire  _GEN_583; // @[LoadQueue.scala 259:25:@9242.4]
  wire  _T_25258; // @[LoadQueue.scala 261:41:@9254.6]
  wire  _GEN_584; // @[LoadQueue.scala 261:62:@9255.6]
  wire  _GEN_585; // @[LoadQueue.scala 259:25:@9250.4]
  wire  _T_25261; // @[LoadQueue.scala 261:41:@9262.6]
  wire  _GEN_586; // @[LoadQueue.scala 261:62:@9263.6]
  wire  _GEN_587; // @[LoadQueue.scala 259:25:@9258.4]
  wire  _T_25264; // @[LoadQueue.scala 261:41:@9270.6]
  wire  _GEN_588; // @[LoadQueue.scala 261:62:@9271.6]
  wire  _GEN_589; // @[LoadQueue.scala 259:25:@9266.4]
  wire  _T_25267; // @[LoadQueue.scala 261:41:@9278.6]
  wire  _GEN_590; // @[LoadQueue.scala 261:62:@9279.6]
  wire  _GEN_591; // @[LoadQueue.scala 259:25:@9274.4]
  wire  _T_25270; // @[LoadQueue.scala 261:41:@9286.6]
  wire  _GEN_592; // @[LoadQueue.scala 261:62:@9287.6]
  wire  _GEN_593; // @[LoadQueue.scala 259:25:@9282.4]
  wire [31:0] _GEN_594; // @[LoadQueue.scala 269:44:@9294.6]
  wire [31:0] _GEN_595; // @[LoadQueue.scala 267:32:@9290.4]
  wire [31:0] _GEN_596; // @[LoadQueue.scala 269:44:@9301.6]
  wire [31:0] _GEN_597; // @[LoadQueue.scala 267:32:@9297.4]
  wire [31:0] _GEN_598; // @[LoadQueue.scala 269:44:@9308.6]
  wire [31:0] _GEN_599; // @[LoadQueue.scala 267:32:@9304.4]
  wire [31:0] _GEN_600; // @[LoadQueue.scala 269:44:@9315.6]
  wire [31:0] _GEN_601; // @[LoadQueue.scala 267:32:@9311.4]
  wire [31:0] _GEN_602; // @[LoadQueue.scala 269:44:@9322.6]
  wire [31:0] _GEN_603; // @[LoadQueue.scala 267:32:@9318.4]
  wire [31:0] _GEN_604; // @[LoadQueue.scala 269:44:@9329.6]
  wire [31:0] _GEN_605; // @[LoadQueue.scala 267:32:@9325.4]
  wire [31:0] _GEN_606; // @[LoadQueue.scala 269:44:@9336.6]
  wire [31:0] _GEN_607; // @[LoadQueue.scala 267:32:@9332.4]
  wire [31:0] _GEN_608; // @[LoadQueue.scala 269:44:@9343.6]
  wire [31:0] _GEN_609; // @[LoadQueue.scala 267:32:@9339.4]
  wire  entriesPorts_0_0; // @[LoadQueue.scala 286:69:@9347.4]
  wire  entriesPorts_0_1; // @[LoadQueue.scala 286:69:@9349.4]
  wire  entriesPorts_0_2; // @[LoadQueue.scala 286:69:@9351.4]
  wire  entriesPorts_0_3; // @[LoadQueue.scala 286:69:@9353.4]
  wire  entriesPorts_0_4; // @[LoadQueue.scala 286:69:@9355.4]
  wire  entriesPorts_0_5; // @[LoadQueue.scala 286:69:@9357.4]
  wire  entriesPorts_0_6; // @[LoadQueue.scala 286:69:@9359.4]
  wire  entriesPorts_0_7; // @[LoadQueue.scala 286:69:@9361.4]
  wire  entriesPorts_1_0; // @[LoadQueue.scala 286:69:@9363.4]
  wire  entriesPorts_1_1; // @[LoadQueue.scala 286:69:@9365.4]
  wire  entriesPorts_1_2; // @[LoadQueue.scala 286:69:@9367.4]
  wire  entriesPorts_1_3; // @[LoadQueue.scala 286:69:@9369.4]
  wire  entriesPorts_1_4; // @[LoadQueue.scala 286:69:@9371.4]
  wire  entriesPorts_1_5; // @[LoadQueue.scala 286:69:@9373.4]
  wire  entriesPorts_1_6; // @[LoadQueue.scala 286:69:@9375.4]
  wire  entriesPorts_1_7; // @[LoadQueue.scala 286:69:@9377.4]
  wire  entriesPorts_2_0; // @[LoadQueue.scala 286:69:@9379.4]
  wire  entriesPorts_2_1; // @[LoadQueue.scala 286:69:@9381.4]
  wire  entriesPorts_2_2; // @[LoadQueue.scala 286:69:@9383.4]
  wire  entriesPorts_2_3; // @[LoadQueue.scala 286:69:@9385.4]
  wire  entriesPorts_2_4; // @[LoadQueue.scala 286:69:@9387.4]
  wire  entriesPorts_2_5; // @[LoadQueue.scala 286:69:@9389.4]
  wire  entriesPorts_2_6; // @[LoadQueue.scala 286:69:@9391.4]
  wire  entriesPorts_2_7; // @[LoadQueue.scala 286:69:@9393.4]
  wire  entriesPorts_3_0; // @[LoadQueue.scala 286:69:@9395.4]
  wire  entriesPorts_3_1; // @[LoadQueue.scala 286:69:@9397.4]
  wire  entriesPorts_3_2; // @[LoadQueue.scala 286:69:@9399.4]
  wire  entriesPorts_3_3; // @[LoadQueue.scala 286:69:@9401.4]
  wire  entriesPorts_3_4; // @[LoadQueue.scala 286:69:@9403.4]
  wire  entriesPorts_3_5; // @[LoadQueue.scala 286:69:@9405.4]
  wire  entriesPorts_3_6; // @[LoadQueue.scala 286:69:@9407.4]
  wire  entriesPorts_3_7; // @[LoadQueue.scala 286:69:@9409.4]
  wire  entriesPorts_4_0; // @[LoadQueue.scala 286:69:@9411.4]
  wire  entriesPorts_4_1; // @[LoadQueue.scala 286:69:@9413.4]
  wire  entriesPorts_4_2; // @[LoadQueue.scala 286:69:@9415.4]
  wire  entriesPorts_4_3; // @[LoadQueue.scala 286:69:@9417.4]
  wire  entriesPorts_4_4; // @[LoadQueue.scala 286:69:@9419.4]
  wire  entriesPorts_4_5; // @[LoadQueue.scala 286:69:@9421.4]
  wire  entriesPorts_4_6; // @[LoadQueue.scala 286:69:@9423.4]
  wire  entriesPorts_4_7; // @[LoadQueue.scala 286:69:@9425.4]
  wire  _T_26091; // @[LoadQueue.scala 298:86:@9429.4]
  wire  _T_26092; // @[LoadQueue.scala 298:83:@9430.4]
  wire  _T_26094; // @[LoadQueue.scala 298:86:@9431.4]
  wire  _T_26095; // @[LoadQueue.scala 298:83:@9432.4]
  wire  _T_26097; // @[LoadQueue.scala 298:86:@9433.4]
  wire  _T_26098; // @[LoadQueue.scala 298:83:@9434.4]
  wire  _T_26100; // @[LoadQueue.scala 298:86:@9435.4]
  wire  _T_26101; // @[LoadQueue.scala 298:83:@9436.4]
  wire  _T_26103; // @[LoadQueue.scala 298:86:@9437.4]
  wire  _T_26104; // @[LoadQueue.scala 298:83:@9438.4]
  wire  _T_26106; // @[LoadQueue.scala 298:86:@9439.4]
  wire  _T_26107; // @[LoadQueue.scala 298:83:@9440.4]
  wire  _T_26109; // @[LoadQueue.scala 298:86:@9441.4]
  wire  _T_26110; // @[LoadQueue.scala 298:83:@9442.4]
  wire  _T_26112; // @[LoadQueue.scala 298:86:@9443.4]
  wire  _T_26113; // @[LoadQueue.scala 298:83:@9444.4]
  wire [7:0] _T_26164; // @[Mux.scala 31:69:@9474.4]
  wire [7:0] _T_26165; // @[Mux.scala 31:69:@9475.4]
  wire [7:0] _T_26166; // @[Mux.scala 31:69:@9476.4]
  wire [7:0] _T_26167; // @[Mux.scala 31:69:@9477.4]
  wire [7:0] _T_26168; // @[Mux.scala 31:69:@9478.4]
  wire [7:0] _T_26169; // @[Mux.scala 31:69:@9479.4]
  wire [7:0] _T_26170; // @[Mux.scala 31:69:@9480.4]
  wire [7:0] _T_26171; // @[Mux.scala 31:69:@9481.4]
  wire  _T_26172; // @[OneHot.scala 66:30:@9482.4]
  wire  _T_26173; // @[OneHot.scala 66:30:@9483.4]
  wire  _T_26174; // @[OneHot.scala 66:30:@9484.4]
  wire  _T_26175; // @[OneHot.scala 66:30:@9485.4]
  wire  _T_26176; // @[OneHot.scala 66:30:@9486.4]
  wire  _T_26177; // @[OneHot.scala 66:30:@9487.4]
  wire  _T_26178; // @[OneHot.scala 66:30:@9488.4]
  wire  _T_26179; // @[OneHot.scala 66:30:@9489.4]
  wire [7:0] _T_26204; // @[Mux.scala 31:69:@9499.4]
  wire [7:0] _T_26205; // @[Mux.scala 31:69:@9500.4]
  wire [7:0] _T_26206; // @[Mux.scala 31:69:@9501.4]
  wire [7:0] _T_26207; // @[Mux.scala 31:69:@9502.4]
  wire [7:0] _T_26208; // @[Mux.scala 31:69:@9503.4]
  wire [7:0] _T_26209; // @[Mux.scala 31:69:@9504.4]
  wire [7:0] _T_26210; // @[Mux.scala 31:69:@9505.4]
  wire [7:0] _T_26211; // @[Mux.scala 31:69:@9506.4]
  wire  _T_26212; // @[OneHot.scala 66:30:@9507.4]
  wire  _T_26213; // @[OneHot.scala 66:30:@9508.4]
  wire  _T_26214; // @[OneHot.scala 66:30:@9509.4]
  wire  _T_26215; // @[OneHot.scala 66:30:@9510.4]
  wire  _T_26216; // @[OneHot.scala 66:30:@9511.4]
  wire  _T_26217; // @[OneHot.scala 66:30:@9512.4]
  wire  _T_26218; // @[OneHot.scala 66:30:@9513.4]
  wire  _T_26219; // @[OneHot.scala 66:30:@9514.4]
  wire [7:0] _T_26244; // @[Mux.scala 31:69:@9524.4]
  wire [7:0] _T_26245; // @[Mux.scala 31:69:@9525.4]
  wire [7:0] _T_26246; // @[Mux.scala 31:69:@9526.4]
  wire [7:0] _T_26247; // @[Mux.scala 31:69:@9527.4]
  wire [7:0] _T_26248; // @[Mux.scala 31:69:@9528.4]
  wire [7:0] _T_26249; // @[Mux.scala 31:69:@9529.4]
  wire [7:0] _T_26250; // @[Mux.scala 31:69:@9530.4]
  wire [7:0] _T_26251; // @[Mux.scala 31:69:@9531.4]
  wire  _T_26252; // @[OneHot.scala 66:30:@9532.4]
  wire  _T_26253; // @[OneHot.scala 66:30:@9533.4]
  wire  _T_26254; // @[OneHot.scala 66:30:@9534.4]
  wire  _T_26255; // @[OneHot.scala 66:30:@9535.4]
  wire  _T_26256; // @[OneHot.scala 66:30:@9536.4]
  wire  _T_26257; // @[OneHot.scala 66:30:@9537.4]
  wire  _T_26258; // @[OneHot.scala 66:30:@9538.4]
  wire  _T_26259; // @[OneHot.scala 66:30:@9539.4]
  wire [7:0] _T_26284; // @[Mux.scala 31:69:@9549.4]
  wire [7:0] _T_26285; // @[Mux.scala 31:69:@9550.4]
  wire [7:0] _T_26286; // @[Mux.scala 31:69:@9551.4]
  wire [7:0] _T_26287; // @[Mux.scala 31:69:@9552.4]
  wire [7:0] _T_26288; // @[Mux.scala 31:69:@9553.4]
  wire [7:0] _T_26289; // @[Mux.scala 31:69:@9554.4]
  wire [7:0] _T_26290; // @[Mux.scala 31:69:@9555.4]
  wire [7:0] _T_26291; // @[Mux.scala 31:69:@9556.4]
  wire  _T_26292; // @[OneHot.scala 66:30:@9557.4]
  wire  _T_26293; // @[OneHot.scala 66:30:@9558.4]
  wire  _T_26294; // @[OneHot.scala 66:30:@9559.4]
  wire  _T_26295; // @[OneHot.scala 66:30:@9560.4]
  wire  _T_26296; // @[OneHot.scala 66:30:@9561.4]
  wire  _T_26297; // @[OneHot.scala 66:30:@9562.4]
  wire  _T_26298; // @[OneHot.scala 66:30:@9563.4]
  wire  _T_26299; // @[OneHot.scala 66:30:@9564.4]
  wire [7:0] _T_26324; // @[Mux.scala 31:69:@9574.4]
  wire [7:0] _T_26325; // @[Mux.scala 31:69:@9575.4]
  wire [7:0] _T_26326; // @[Mux.scala 31:69:@9576.4]
  wire [7:0] _T_26327; // @[Mux.scala 31:69:@9577.4]
  wire [7:0] _T_26328; // @[Mux.scala 31:69:@9578.4]
  wire [7:0] _T_26329; // @[Mux.scala 31:69:@9579.4]
  wire [7:0] _T_26330; // @[Mux.scala 31:69:@9580.4]
  wire [7:0] _T_26331; // @[Mux.scala 31:69:@9581.4]
  wire  _T_26332; // @[OneHot.scala 66:30:@9582.4]
  wire  _T_26333; // @[OneHot.scala 66:30:@9583.4]
  wire  _T_26334; // @[OneHot.scala 66:30:@9584.4]
  wire  _T_26335; // @[OneHot.scala 66:30:@9585.4]
  wire  _T_26336; // @[OneHot.scala 66:30:@9586.4]
  wire  _T_26337; // @[OneHot.scala 66:30:@9587.4]
  wire  _T_26338; // @[OneHot.scala 66:30:@9588.4]
  wire  _T_26339; // @[OneHot.scala 66:30:@9589.4]
  wire [7:0] _T_26364; // @[Mux.scala 31:69:@9599.4]
  wire [7:0] _T_26365; // @[Mux.scala 31:69:@9600.4]
  wire [7:0] _T_26366; // @[Mux.scala 31:69:@9601.4]
  wire [7:0] _T_26367; // @[Mux.scala 31:69:@9602.4]
  wire [7:0] _T_26368; // @[Mux.scala 31:69:@9603.4]
  wire [7:0] _T_26369; // @[Mux.scala 31:69:@9604.4]
  wire [7:0] _T_26370; // @[Mux.scala 31:69:@9605.4]
  wire [7:0] _T_26371; // @[Mux.scala 31:69:@9606.4]
  wire  _T_26372; // @[OneHot.scala 66:30:@9607.4]
  wire  _T_26373; // @[OneHot.scala 66:30:@9608.4]
  wire  _T_26374; // @[OneHot.scala 66:30:@9609.4]
  wire  _T_26375; // @[OneHot.scala 66:30:@9610.4]
  wire  _T_26376; // @[OneHot.scala 66:30:@9611.4]
  wire  _T_26377; // @[OneHot.scala 66:30:@9612.4]
  wire  _T_26378; // @[OneHot.scala 66:30:@9613.4]
  wire  _T_26379; // @[OneHot.scala 66:30:@9614.4]
  wire [7:0] _T_26404; // @[Mux.scala 31:69:@9624.4]
  wire [7:0] _T_26405; // @[Mux.scala 31:69:@9625.4]
  wire [7:0] _T_26406; // @[Mux.scala 31:69:@9626.4]
  wire [7:0] _T_26407; // @[Mux.scala 31:69:@9627.4]
  wire [7:0] _T_26408; // @[Mux.scala 31:69:@9628.4]
  wire [7:0] _T_26409; // @[Mux.scala 31:69:@9629.4]
  wire [7:0] _T_26410; // @[Mux.scala 31:69:@9630.4]
  wire [7:0] _T_26411; // @[Mux.scala 31:69:@9631.4]
  wire  _T_26412; // @[OneHot.scala 66:30:@9632.4]
  wire  _T_26413; // @[OneHot.scala 66:30:@9633.4]
  wire  _T_26414; // @[OneHot.scala 66:30:@9634.4]
  wire  _T_26415; // @[OneHot.scala 66:30:@9635.4]
  wire  _T_26416; // @[OneHot.scala 66:30:@9636.4]
  wire  _T_26417; // @[OneHot.scala 66:30:@9637.4]
  wire  _T_26418; // @[OneHot.scala 66:30:@9638.4]
  wire  _T_26419; // @[OneHot.scala 66:30:@9639.4]
  wire [7:0] _T_26444; // @[Mux.scala 31:69:@9649.4]
  wire [7:0] _T_26445; // @[Mux.scala 31:69:@9650.4]
  wire [7:0] _T_26446; // @[Mux.scala 31:69:@9651.4]
  wire [7:0] _T_26447; // @[Mux.scala 31:69:@9652.4]
  wire [7:0] _T_26448; // @[Mux.scala 31:69:@9653.4]
  wire [7:0] _T_26449; // @[Mux.scala 31:69:@9654.4]
  wire [7:0] _T_26450; // @[Mux.scala 31:69:@9655.4]
  wire [7:0] _T_26451; // @[Mux.scala 31:69:@9656.4]
  wire  _T_26452; // @[OneHot.scala 66:30:@9657.4]
  wire  _T_26453; // @[OneHot.scala 66:30:@9658.4]
  wire  _T_26454; // @[OneHot.scala 66:30:@9659.4]
  wire  _T_26455; // @[OneHot.scala 66:30:@9660.4]
  wire  _T_26456; // @[OneHot.scala 66:30:@9661.4]
  wire  _T_26457; // @[OneHot.scala 66:30:@9662.4]
  wire  _T_26458; // @[OneHot.scala 66:30:@9663.4]
  wire  _T_26459; // @[OneHot.scala 66:30:@9664.4]
  wire [7:0] _T_26500; // @[Mux.scala 19:72:@9680.4]
  wire [7:0] _T_26502; // @[Mux.scala 19:72:@9681.4]
  wire [7:0] _T_26509; // @[Mux.scala 19:72:@9688.4]
  wire [7:0] _T_26511; // @[Mux.scala 19:72:@9689.4]
  wire [7:0] _T_26518; // @[Mux.scala 19:72:@9696.4]
  wire [7:0] _T_26520; // @[Mux.scala 19:72:@9697.4]
  wire [7:0] _T_26527; // @[Mux.scala 19:72:@9704.4]
  wire [7:0] _T_26529; // @[Mux.scala 19:72:@9705.4]
  wire [7:0] _T_26536; // @[Mux.scala 19:72:@9712.4]
  wire [7:0] _T_26538; // @[Mux.scala 19:72:@9713.4]
  wire [7:0] _T_26545; // @[Mux.scala 19:72:@9720.4]
  wire [7:0] _T_26547; // @[Mux.scala 19:72:@9721.4]
  wire [7:0] _T_26554; // @[Mux.scala 19:72:@9728.4]
  wire [7:0] _T_26556; // @[Mux.scala 19:72:@9729.4]
  wire [7:0] _T_26563; // @[Mux.scala 19:72:@9736.4]
  wire [7:0] _T_26565; // @[Mux.scala 19:72:@9737.4]
  wire [7:0] _T_26566; // @[Mux.scala 19:72:@9738.4]
  wire [7:0] _T_26567; // @[Mux.scala 19:72:@9739.4]
  wire [7:0] _T_26568; // @[Mux.scala 19:72:@9740.4]
  wire [7:0] _T_26569; // @[Mux.scala 19:72:@9741.4]
  wire [7:0] _T_26570; // @[Mux.scala 19:72:@9742.4]
  wire [7:0] _T_26571; // @[Mux.scala 19:72:@9743.4]
  wire [7:0] _T_26572; // @[Mux.scala 19:72:@9744.4]
  wire  inputPriorityPorts_0_0; // @[Mux.scala 19:72:@9748.4]
  wire  inputPriorityPorts_0_1; // @[Mux.scala 19:72:@9750.4]
  wire  inputPriorityPorts_0_2; // @[Mux.scala 19:72:@9752.4]
  wire  inputPriorityPorts_0_3; // @[Mux.scala 19:72:@9754.4]
  wire  inputPriorityPorts_0_4; // @[Mux.scala 19:72:@9756.4]
  wire  inputPriorityPorts_0_5; // @[Mux.scala 19:72:@9758.4]
  wire  inputPriorityPorts_0_6; // @[Mux.scala 19:72:@9760.4]
  wire  inputPriorityPorts_0_7; // @[Mux.scala 19:72:@9762.4]
  wire [7:0] _T_26686; // @[Mux.scala 31:69:@9792.4]
  wire [7:0] _T_26687; // @[Mux.scala 31:69:@9793.4]
  wire [7:0] _T_26688; // @[Mux.scala 31:69:@9794.4]
  wire [7:0] _T_26689; // @[Mux.scala 31:69:@9795.4]
  wire [7:0] _T_26690; // @[Mux.scala 31:69:@9796.4]
  wire [7:0] _T_26691; // @[Mux.scala 31:69:@9797.4]
  wire [7:0] _T_26692; // @[Mux.scala 31:69:@9798.4]
  wire [7:0] _T_26693; // @[Mux.scala 31:69:@9799.4]
  wire  _T_26694; // @[OneHot.scala 66:30:@9800.4]
  wire  _T_26695; // @[OneHot.scala 66:30:@9801.4]
  wire  _T_26696; // @[OneHot.scala 66:30:@9802.4]
  wire  _T_26697; // @[OneHot.scala 66:30:@9803.4]
  wire  _T_26698; // @[OneHot.scala 66:30:@9804.4]
  wire  _T_26699; // @[OneHot.scala 66:30:@9805.4]
  wire  _T_26700; // @[OneHot.scala 66:30:@9806.4]
  wire  _T_26701; // @[OneHot.scala 66:30:@9807.4]
  wire [7:0] _T_26726; // @[Mux.scala 31:69:@9817.4]
  wire [7:0] _T_26727; // @[Mux.scala 31:69:@9818.4]
  wire [7:0] _T_26728; // @[Mux.scala 31:69:@9819.4]
  wire [7:0] _T_26729; // @[Mux.scala 31:69:@9820.4]
  wire [7:0] _T_26730; // @[Mux.scala 31:69:@9821.4]
  wire [7:0] _T_26731; // @[Mux.scala 31:69:@9822.4]
  wire [7:0] _T_26732; // @[Mux.scala 31:69:@9823.4]
  wire [7:0] _T_26733; // @[Mux.scala 31:69:@9824.4]
  wire  _T_26734; // @[OneHot.scala 66:30:@9825.4]
  wire  _T_26735; // @[OneHot.scala 66:30:@9826.4]
  wire  _T_26736; // @[OneHot.scala 66:30:@9827.4]
  wire  _T_26737; // @[OneHot.scala 66:30:@9828.4]
  wire  _T_26738; // @[OneHot.scala 66:30:@9829.4]
  wire  _T_26739; // @[OneHot.scala 66:30:@9830.4]
  wire  _T_26740; // @[OneHot.scala 66:30:@9831.4]
  wire  _T_26741; // @[OneHot.scala 66:30:@9832.4]
  wire [7:0] _T_26766; // @[Mux.scala 31:69:@9842.4]
  wire [7:0] _T_26767; // @[Mux.scala 31:69:@9843.4]
  wire [7:0] _T_26768; // @[Mux.scala 31:69:@9844.4]
  wire [7:0] _T_26769; // @[Mux.scala 31:69:@9845.4]
  wire [7:0] _T_26770; // @[Mux.scala 31:69:@9846.4]
  wire [7:0] _T_26771; // @[Mux.scala 31:69:@9847.4]
  wire [7:0] _T_26772; // @[Mux.scala 31:69:@9848.4]
  wire [7:0] _T_26773; // @[Mux.scala 31:69:@9849.4]
  wire  _T_26774; // @[OneHot.scala 66:30:@9850.4]
  wire  _T_26775; // @[OneHot.scala 66:30:@9851.4]
  wire  _T_26776; // @[OneHot.scala 66:30:@9852.4]
  wire  _T_26777; // @[OneHot.scala 66:30:@9853.4]
  wire  _T_26778; // @[OneHot.scala 66:30:@9854.4]
  wire  _T_26779; // @[OneHot.scala 66:30:@9855.4]
  wire  _T_26780; // @[OneHot.scala 66:30:@9856.4]
  wire  _T_26781; // @[OneHot.scala 66:30:@9857.4]
  wire [7:0] _T_26806; // @[Mux.scala 31:69:@9867.4]
  wire [7:0] _T_26807; // @[Mux.scala 31:69:@9868.4]
  wire [7:0] _T_26808; // @[Mux.scala 31:69:@9869.4]
  wire [7:0] _T_26809; // @[Mux.scala 31:69:@9870.4]
  wire [7:0] _T_26810; // @[Mux.scala 31:69:@9871.4]
  wire [7:0] _T_26811; // @[Mux.scala 31:69:@9872.4]
  wire [7:0] _T_26812; // @[Mux.scala 31:69:@9873.4]
  wire [7:0] _T_26813; // @[Mux.scala 31:69:@9874.4]
  wire  _T_26814; // @[OneHot.scala 66:30:@9875.4]
  wire  _T_26815; // @[OneHot.scala 66:30:@9876.4]
  wire  _T_26816; // @[OneHot.scala 66:30:@9877.4]
  wire  _T_26817; // @[OneHot.scala 66:30:@9878.4]
  wire  _T_26818; // @[OneHot.scala 66:30:@9879.4]
  wire  _T_26819; // @[OneHot.scala 66:30:@9880.4]
  wire  _T_26820; // @[OneHot.scala 66:30:@9881.4]
  wire  _T_26821; // @[OneHot.scala 66:30:@9882.4]
  wire [7:0] _T_26846; // @[Mux.scala 31:69:@9892.4]
  wire [7:0] _T_26847; // @[Mux.scala 31:69:@9893.4]
  wire [7:0] _T_26848; // @[Mux.scala 31:69:@9894.4]
  wire [7:0] _T_26849; // @[Mux.scala 31:69:@9895.4]
  wire [7:0] _T_26850; // @[Mux.scala 31:69:@9896.4]
  wire [7:0] _T_26851; // @[Mux.scala 31:69:@9897.4]
  wire [7:0] _T_26852; // @[Mux.scala 31:69:@9898.4]
  wire [7:0] _T_26853; // @[Mux.scala 31:69:@9899.4]
  wire  _T_26854; // @[OneHot.scala 66:30:@9900.4]
  wire  _T_26855; // @[OneHot.scala 66:30:@9901.4]
  wire  _T_26856; // @[OneHot.scala 66:30:@9902.4]
  wire  _T_26857; // @[OneHot.scala 66:30:@9903.4]
  wire  _T_26858; // @[OneHot.scala 66:30:@9904.4]
  wire  _T_26859; // @[OneHot.scala 66:30:@9905.4]
  wire  _T_26860; // @[OneHot.scala 66:30:@9906.4]
  wire  _T_26861; // @[OneHot.scala 66:30:@9907.4]
  wire [7:0] _T_26886; // @[Mux.scala 31:69:@9917.4]
  wire [7:0] _T_26887; // @[Mux.scala 31:69:@9918.4]
  wire [7:0] _T_26888; // @[Mux.scala 31:69:@9919.4]
  wire [7:0] _T_26889; // @[Mux.scala 31:69:@9920.4]
  wire [7:0] _T_26890; // @[Mux.scala 31:69:@9921.4]
  wire [7:0] _T_26891; // @[Mux.scala 31:69:@9922.4]
  wire [7:0] _T_26892; // @[Mux.scala 31:69:@9923.4]
  wire [7:0] _T_26893; // @[Mux.scala 31:69:@9924.4]
  wire  _T_26894; // @[OneHot.scala 66:30:@9925.4]
  wire  _T_26895; // @[OneHot.scala 66:30:@9926.4]
  wire  _T_26896; // @[OneHot.scala 66:30:@9927.4]
  wire  _T_26897; // @[OneHot.scala 66:30:@9928.4]
  wire  _T_26898; // @[OneHot.scala 66:30:@9929.4]
  wire  _T_26899; // @[OneHot.scala 66:30:@9930.4]
  wire  _T_26900; // @[OneHot.scala 66:30:@9931.4]
  wire  _T_26901; // @[OneHot.scala 66:30:@9932.4]
  wire [7:0] _T_26926; // @[Mux.scala 31:69:@9942.4]
  wire [7:0] _T_26927; // @[Mux.scala 31:69:@9943.4]
  wire [7:0] _T_26928; // @[Mux.scala 31:69:@9944.4]
  wire [7:0] _T_26929; // @[Mux.scala 31:69:@9945.4]
  wire [7:0] _T_26930; // @[Mux.scala 31:69:@9946.4]
  wire [7:0] _T_26931; // @[Mux.scala 31:69:@9947.4]
  wire [7:0] _T_26932; // @[Mux.scala 31:69:@9948.4]
  wire [7:0] _T_26933; // @[Mux.scala 31:69:@9949.4]
  wire  _T_26934; // @[OneHot.scala 66:30:@9950.4]
  wire  _T_26935; // @[OneHot.scala 66:30:@9951.4]
  wire  _T_26936; // @[OneHot.scala 66:30:@9952.4]
  wire  _T_26937; // @[OneHot.scala 66:30:@9953.4]
  wire  _T_26938; // @[OneHot.scala 66:30:@9954.4]
  wire  _T_26939; // @[OneHot.scala 66:30:@9955.4]
  wire  _T_26940; // @[OneHot.scala 66:30:@9956.4]
  wire  _T_26941; // @[OneHot.scala 66:30:@9957.4]
  wire [7:0] _T_26966; // @[Mux.scala 31:69:@9967.4]
  wire [7:0] _T_26967; // @[Mux.scala 31:69:@9968.4]
  wire [7:0] _T_26968; // @[Mux.scala 31:69:@9969.4]
  wire [7:0] _T_26969; // @[Mux.scala 31:69:@9970.4]
  wire [7:0] _T_26970; // @[Mux.scala 31:69:@9971.4]
  wire [7:0] _T_26971; // @[Mux.scala 31:69:@9972.4]
  wire [7:0] _T_26972; // @[Mux.scala 31:69:@9973.4]
  wire [7:0] _T_26973; // @[Mux.scala 31:69:@9974.4]
  wire  _T_26974; // @[OneHot.scala 66:30:@9975.4]
  wire  _T_26975; // @[OneHot.scala 66:30:@9976.4]
  wire  _T_26976; // @[OneHot.scala 66:30:@9977.4]
  wire  _T_26977; // @[OneHot.scala 66:30:@9978.4]
  wire  _T_26978; // @[OneHot.scala 66:30:@9979.4]
  wire  _T_26979; // @[OneHot.scala 66:30:@9980.4]
  wire  _T_26980; // @[OneHot.scala 66:30:@9981.4]
  wire  _T_26981; // @[OneHot.scala 66:30:@9982.4]
  wire [7:0] _T_27022; // @[Mux.scala 19:72:@9998.4]
  wire [7:0] _T_27024; // @[Mux.scala 19:72:@9999.4]
  wire [7:0] _T_27031; // @[Mux.scala 19:72:@10006.4]
  wire [7:0] _T_27033; // @[Mux.scala 19:72:@10007.4]
  wire [7:0] _T_27040; // @[Mux.scala 19:72:@10014.4]
  wire [7:0] _T_27042; // @[Mux.scala 19:72:@10015.4]
  wire [7:0] _T_27049; // @[Mux.scala 19:72:@10022.4]
  wire [7:0] _T_27051; // @[Mux.scala 19:72:@10023.4]
  wire [7:0] _T_27058; // @[Mux.scala 19:72:@10030.4]
  wire [7:0] _T_27060; // @[Mux.scala 19:72:@10031.4]
  wire [7:0] _T_27067; // @[Mux.scala 19:72:@10038.4]
  wire [7:0] _T_27069; // @[Mux.scala 19:72:@10039.4]
  wire [7:0] _T_27076; // @[Mux.scala 19:72:@10046.4]
  wire [7:0] _T_27078; // @[Mux.scala 19:72:@10047.4]
  wire [7:0] _T_27085; // @[Mux.scala 19:72:@10054.4]
  wire [7:0] _T_27087; // @[Mux.scala 19:72:@10055.4]
  wire [7:0] _T_27088; // @[Mux.scala 19:72:@10056.4]
  wire [7:0] _T_27089; // @[Mux.scala 19:72:@10057.4]
  wire [7:0] _T_27090; // @[Mux.scala 19:72:@10058.4]
  wire [7:0] _T_27091; // @[Mux.scala 19:72:@10059.4]
  wire [7:0] _T_27092; // @[Mux.scala 19:72:@10060.4]
  wire [7:0] _T_27093; // @[Mux.scala 19:72:@10061.4]
  wire [7:0] _T_27094; // @[Mux.scala 19:72:@10062.4]
  wire  outputPriorityPorts_0_0; // @[Mux.scala 19:72:@10066.4]
  wire  outputPriorityPorts_0_1; // @[Mux.scala 19:72:@10068.4]
  wire  outputPriorityPorts_0_2; // @[Mux.scala 19:72:@10070.4]
  wire  outputPriorityPorts_0_3; // @[Mux.scala 19:72:@10072.4]
  wire  outputPriorityPorts_0_4; // @[Mux.scala 19:72:@10074.4]
  wire  outputPriorityPorts_0_5; // @[Mux.scala 19:72:@10076.4]
  wire  outputPriorityPorts_0_6; // @[Mux.scala 19:72:@10078.4]
  wire  outputPriorityPorts_0_7; // @[Mux.scala 19:72:@10080.4]
  wire  _T_27174; // @[LoadQueue.scala 298:83:@10091.4]
  wire  _T_27177; // @[LoadQueue.scala 298:83:@10093.4]
  wire  _T_27180; // @[LoadQueue.scala 298:83:@10095.4]
  wire  _T_27183; // @[LoadQueue.scala 298:83:@10097.4]
  wire  _T_27186; // @[LoadQueue.scala 298:83:@10099.4]
  wire  _T_27189; // @[LoadQueue.scala 298:83:@10101.4]
  wire  _T_27192; // @[LoadQueue.scala 298:83:@10103.4]
  wire  _T_27195; // @[LoadQueue.scala 298:83:@10105.4]
  wire [7:0] _T_27246; // @[Mux.scala 31:69:@10135.4]
  wire [7:0] _T_27247; // @[Mux.scala 31:69:@10136.4]
  wire [7:0] _T_27248; // @[Mux.scala 31:69:@10137.4]
  wire [7:0] _T_27249; // @[Mux.scala 31:69:@10138.4]
  wire [7:0] _T_27250; // @[Mux.scala 31:69:@10139.4]
  wire [7:0] _T_27251; // @[Mux.scala 31:69:@10140.4]
  wire [7:0] _T_27252; // @[Mux.scala 31:69:@10141.4]
  wire [7:0] _T_27253; // @[Mux.scala 31:69:@10142.4]
  wire  _T_27254; // @[OneHot.scala 66:30:@10143.4]
  wire  _T_27255; // @[OneHot.scala 66:30:@10144.4]
  wire  _T_27256; // @[OneHot.scala 66:30:@10145.4]
  wire  _T_27257; // @[OneHot.scala 66:30:@10146.4]
  wire  _T_27258; // @[OneHot.scala 66:30:@10147.4]
  wire  _T_27259; // @[OneHot.scala 66:30:@10148.4]
  wire  _T_27260; // @[OneHot.scala 66:30:@10149.4]
  wire  _T_27261; // @[OneHot.scala 66:30:@10150.4]
  wire [7:0] _T_27286; // @[Mux.scala 31:69:@10160.4]
  wire [7:0] _T_27287; // @[Mux.scala 31:69:@10161.4]
  wire [7:0] _T_27288; // @[Mux.scala 31:69:@10162.4]
  wire [7:0] _T_27289; // @[Mux.scala 31:69:@10163.4]
  wire [7:0] _T_27290; // @[Mux.scala 31:69:@10164.4]
  wire [7:0] _T_27291; // @[Mux.scala 31:69:@10165.4]
  wire [7:0] _T_27292; // @[Mux.scala 31:69:@10166.4]
  wire [7:0] _T_27293; // @[Mux.scala 31:69:@10167.4]
  wire  _T_27294; // @[OneHot.scala 66:30:@10168.4]
  wire  _T_27295; // @[OneHot.scala 66:30:@10169.4]
  wire  _T_27296; // @[OneHot.scala 66:30:@10170.4]
  wire  _T_27297; // @[OneHot.scala 66:30:@10171.4]
  wire  _T_27298; // @[OneHot.scala 66:30:@10172.4]
  wire  _T_27299; // @[OneHot.scala 66:30:@10173.4]
  wire  _T_27300; // @[OneHot.scala 66:30:@10174.4]
  wire  _T_27301; // @[OneHot.scala 66:30:@10175.4]
  wire [7:0] _T_27326; // @[Mux.scala 31:69:@10185.4]
  wire [7:0] _T_27327; // @[Mux.scala 31:69:@10186.4]
  wire [7:0] _T_27328; // @[Mux.scala 31:69:@10187.4]
  wire [7:0] _T_27329; // @[Mux.scala 31:69:@10188.4]
  wire [7:0] _T_27330; // @[Mux.scala 31:69:@10189.4]
  wire [7:0] _T_27331; // @[Mux.scala 31:69:@10190.4]
  wire [7:0] _T_27332; // @[Mux.scala 31:69:@10191.4]
  wire [7:0] _T_27333; // @[Mux.scala 31:69:@10192.4]
  wire  _T_27334; // @[OneHot.scala 66:30:@10193.4]
  wire  _T_27335; // @[OneHot.scala 66:30:@10194.4]
  wire  _T_27336; // @[OneHot.scala 66:30:@10195.4]
  wire  _T_27337; // @[OneHot.scala 66:30:@10196.4]
  wire  _T_27338; // @[OneHot.scala 66:30:@10197.4]
  wire  _T_27339; // @[OneHot.scala 66:30:@10198.4]
  wire  _T_27340; // @[OneHot.scala 66:30:@10199.4]
  wire  _T_27341; // @[OneHot.scala 66:30:@10200.4]
  wire [7:0] _T_27366; // @[Mux.scala 31:69:@10210.4]
  wire [7:0] _T_27367; // @[Mux.scala 31:69:@10211.4]
  wire [7:0] _T_27368; // @[Mux.scala 31:69:@10212.4]
  wire [7:0] _T_27369; // @[Mux.scala 31:69:@10213.4]
  wire [7:0] _T_27370; // @[Mux.scala 31:69:@10214.4]
  wire [7:0] _T_27371; // @[Mux.scala 31:69:@10215.4]
  wire [7:0] _T_27372; // @[Mux.scala 31:69:@10216.4]
  wire [7:0] _T_27373; // @[Mux.scala 31:69:@10217.4]
  wire  _T_27374; // @[OneHot.scala 66:30:@10218.4]
  wire  _T_27375; // @[OneHot.scala 66:30:@10219.4]
  wire  _T_27376; // @[OneHot.scala 66:30:@10220.4]
  wire  _T_27377; // @[OneHot.scala 66:30:@10221.4]
  wire  _T_27378; // @[OneHot.scala 66:30:@10222.4]
  wire  _T_27379; // @[OneHot.scala 66:30:@10223.4]
  wire  _T_27380; // @[OneHot.scala 66:30:@10224.4]
  wire  _T_27381; // @[OneHot.scala 66:30:@10225.4]
  wire [7:0] _T_27406; // @[Mux.scala 31:69:@10235.4]
  wire [7:0] _T_27407; // @[Mux.scala 31:69:@10236.4]
  wire [7:0] _T_27408; // @[Mux.scala 31:69:@10237.4]
  wire [7:0] _T_27409; // @[Mux.scala 31:69:@10238.4]
  wire [7:0] _T_27410; // @[Mux.scala 31:69:@10239.4]
  wire [7:0] _T_27411; // @[Mux.scala 31:69:@10240.4]
  wire [7:0] _T_27412; // @[Mux.scala 31:69:@10241.4]
  wire [7:0] _T_27413; // @[Mux.scala 31:69:@10242.4]
  wire  _T_27414; // @[OneHot.scala 66:30:@10243.4]
  wire  _T_27415; // @[OneHot.scala 66:30:@10244.4]
  wire  _T_27416; // @[OneHot.scala 66:30:@10245.4]
  wire  _T_27417; // @[OneHot.scala 66:30:@10246.4]
  wire  _T_27418; // @[OneHot.scala 66:30:@10247.4]
  wire  _T_27419; // @[OneHot.scala 66:30:@10248.4]
  wire  _T_27420; // @[OneHot.scala 66:30:@10249.4]
  wire  _T_27421; // @[OneHot.scala 66:30:@10250.4]
  wire [7:0] _T_27446; // @[Mux.scala 31:69:@10260.4]
  wire [7:0] _T_27447; // @[Mux.scala 31:69:@10261.4]
  wire [7:0] _T_27448; // @[Mux.scala 31:69:@10262.4]
  wire [7:0] _T_27449; // @[Mux.scala 31:69:@10263.4]
  wire [7:0] _T_27450; // @[Mux.scala 31:69:@10264.4]
  wire [7:0] _T_27451; // @[Mux.scala 31:69:@10265.4]
  wire [7:0] _T_27452; // @[Mux.scala 31:69:@10266.4]
  wire [7:0] _T_27453; // @[Mux.scala 31:69:@10267.4]
  wire  _T_27454; // @[OneHot.scala 66:30:@10268.4]
  wire  _T_27455; // @[OneHot.scala 66:30:@10269.4]
  wire  _T_27456; // @[OneHot.scala 66:30:@10270.4]
  wire  _T_27457; // @[OneHot.scala 66:30:@10271.4]
  wire  _T_27458; // @[OneHot.scala 66:30:@10272.4]
  wire  _T_27459; // @[OneHot.scala 66:30:@10273.4]
  wire  _T_27460; // @[OneHot.scala 66:30:@10274.4]
  wire  _T_27461; // @[OneHot.scala 66:30:@10275.4]
  wire [7:0] _T_27486; // @[Mux.scala 31:69:@10285.4]
  wire [7:0] _T_27487; // @[Mux.scala 31:69:@10286.4]
  wire [7:0] _T_27488; // @[Mux.scala 31:69:@10287.4]
  wire [7:0] _T_27489; // @[Mux.scala 31:69:@10288.4]
  wire [7:0] _T_27490; // @[Mux.scala 31:69:@10289.4]
  wire [7:0] _T_27491; // @[Mux.scala 31:69:@10290.4]
  wire [7:0] _T_27492; // @[Mux.scala 31:69:@10291.4]
  wire [7:0] _T_27493; // @[Mux.scala 31:69:@10292.4]
  wire  _T_27494; // @[OneHot.scala 66:30:@10293.4]
  wire  _T_27495; // @[OneHot.scala 66:30:@10294.4]
  wire  _T_27496; // @[OneHot.scala 66:30:@10295.4]
  wire  _T_27497; // @[OneHot.scala 66:30:@10296.4]
  wire  _T_27498; // @[OneHot.scala 66:30:@10297.4]
  wire  _T_27499; // @[OneHot.scala 66:30:@10298.4]
  wire  _T_27500; // @[OneHot.scala 66:30:@10299.4]
  wire  _T_27501; // @[OneHot.scala 66:30:@10300.4]
  wire [7:0] _T_27526; // @[Mux.scala 31:69:@10310.4]
  wire [7:0] _T_27527; // @[Mux.scala 31:69:@10311.4]
  wire [7:0] _T_27528; // @[Mux.scala 31:69:@10312.4]
  wire [7:0] _T_27529; // @[Mux.scala 31:69:@10313.4]
  wire [7:0] _T_27530; // @[Mux.scala 31:69:@10314.4]
  wire [7:0] _T_27531; // @[Mux.scala 31:69:@10315.4]
  wire [7:0] _T_27532; // @[Mux.scala 31:69:@10316.4]
  wire [7:0] _T_27533; // @[Mux.scala 31:69:@10317.4]
  wire  _T_27534; // @[OneHot.scala 66:30:@10318.4]
  wire  _T_27535; // @[OneHot.scala 66:30:@10319.4]
  wire  _T_27536; // @[OneHot.scala 66:30:@10320.4]
  wire  _T_27537; // @[OneHot.scala 66:30:@10321.4]
  wire  _T_27538; // @[OneHot.scala 66:30:@10322.4]
  wire  _T_27539; // @[OneHot.scala 66:30:@10323.4]
  wire  _T_27540; // @[OneHot.scala 66:30:@10324.4]
  wire  _T_27541; // @[OneHot.scala 66:30:@10325.4]
  wire [7:0] _T_27582; // @[Mux.scala 19:72:@10341.4]
  wire [7:0] _T_27584; // @[Mux.scala 19:72:@10342.4]
  wire [7:0] _T_27591; // @[Mux.scala 19:72:@10349.4]
  wire [7:0] _T_27593; // @[Mux.scala 19:72:@10350.4]
  wire [7:0] _T_27600; // @[Mux.scala 19:72:@10357.4]
  wire [7:0] _T_27602; // @[Mux.scala 19:72:@10358.4]
  wire [7:0] _T_27609; // @[Mux.scala 19:72:@10365.4]
  wire [7:0] _T_27611; // @[Mux.scala 19:72:@10366.4]
  wire [7:0] _T_27618; // @[Mux.scala 19:72:@10373.4]
  wire [7:0] _T_27620; // @[Mux.scala 19:72:@10374.4]
  wire [7:0] _T_27627; // @[Mux.scala 19:72:@10381.4]
  wire [7:0] _T_27629; // @[Mux.scala 19:72:@10382.4]
  wire [7:0] _T_27636; // @[Mux.scala 19:72:@10389.4]
  wire [7:0] _T_27638; // @[Mux.scala 19:72:@10390.4]
  wire [7:0] _T_27645; // @[Mux.scala 19:72:@10397.4]
  wire [7:0] _T_27647; // @[Mux.scala 19:72:@10398.4]
  wire [7:0] _T_27648; // @[Mux.scala 19:72:@10399.4]
  wire [7:0] _T_27649; // @[Mux.scala 19:72:@10400.4]
  wire [7:0] _T_27650; // @[Mux.scala 19:72:@10401.4]
  wire [7:0] _T_27651; // @[Mux.scala 19:72:@10402.4]
  wire [7:0] _T_27652; // @[Mux.scala 19:72:@10403.4]
  wire [7:0] _T_27653; // @[Mux.scala 19:72:@10404.4]
  wire [7:0] _T_27654; // @[Mux.scala 19:72:@10405.4]
  wire  inputPriorityPorts_1_0; // @[Mux.scala 19:72:@10409.4]
  wire  inputPriorityPorts_1_1; // @[Mux.scala 19:72:@10411.4]
  wire  inputPriorityPorts_1_2; // @[Mux.scala 19:72:@10413.4]
  wire  inputPriorityPorts_1_3; // @[Mux.scala 19:72:@10415.4]
  wire  inputPriorityPorts_1_4; // @[Mux.scala 19:72:@10417.4]
  wire  inputPriorityPorts_1_5; // @[Mux.scala 19:72:@10419.4]
  wire  inputPriorityPorts_1_6; // @[Mux.scala 19:72:@10421.4]
  wire  inputPriorityPorts_1_7; // @[Mux.scala 19:72:@10423.4]
  wire [7:0] _T_27768; // @[Mux.scala 31:69:@10453.4]
  wire [7:0] _T_27769; // @[Mux.scala 31:69:@10454.4]
  wire [7:0] _T_27770; // @[Mux.scala 31:69:@10455.4]
  wire [7:0] _T_27771; // @[Mux.scala 31:69:@10456.4]
  wire [7:0] _T_27772; // @[Mux.scala 31:69:@10457.4]
  wire [7:0] _T_27773; // @[Mux.scala 31:69:@10458.4]
  wire [7:0] _T_27774; // @[Mux.scala 31:69:@10459.4]
  wire [7:0] _T_27775; // @[Mux.scala 31:69:@10460.4]
  wire  _T_27776; // @[OneHot.scala 66:30:@10461.4]
  wire  _T_27777; // @[OneHot.scala 66:30:@10462.4]
  wire  _T_27778; // @[OneHot.scala 66:30:@10463.4]
  wire  _T_27779; // @[OneHot.scala 66:30:@10464.4]
  wire  _T_27780; // @[OneHot.scala 66:30:@10465.4]
  wire  _T_27781; // @[OneHot.scala 66:30:@10466.4]
  wire  _T_27782; // @[OneHot.scala 66:30:@10467.4]
  wire  _T_27783; // @[OneHot.scala 66:30:@10468.4]
  wire [7:0] _T_27808; // @[Mux.scala 31:69:@10478.4]
  wire [7:0] _T_27809; // @[Mux.scala 31:69:@10479.4]
  wire [7:0] _T_27810; // @[Mux.scala 31:69:@10480.4]
  wire [7:0] _T_27811; // @[Mux.scala 31:69:@10481.4]
  wire [7:0] _T_27812; // @[Mux.scala 31:69:@10482.4]
  wire [7:0] _T_27813; // @[Mux.scala 31:69:@10483.4]
  wire [7:0] _T_27814; // @[Mux.scala 31:69:@10484.4]
  wire [7:0] _T_27815; // @[Mux.scala 31:69:@10485.4]
  wire  _T_27816; // @[OneHot.scala 66:30:@10486.4]
  wire  _T_27817; // @[OneHot.scala 66:30:@10487.4]
  wire  _T_27818; // @[OneHot.scala 66:30:@10488.4]
  wire  _T_27819; // @[OneHot.scala 66:30:@10489.4]
  wire  _T_27820; // @[OneHot.scala 66:30:@10490.4]
  wire  _T_27821; // @[OneHot.scala 66:30:@10491.4]
  wire  _T_27822; // @[OneHot.scala 66:30:@10492.4]
  wire  _T_27823; // @[OneHot.scala 66:30:@10493.4]
  wire [7:0] _T_27848; // @[Mux.scala 31:69:@10503.4]
  wire [7:0] _T_27849; // @[Mux.scala 31:69:@10504.4]
  wire [7:0] _T_27850; // @[Mux.scala 31:69:@10505.4]
  wire [7:0] _T_27851; // @[Mux.scala 31:69:@10506.4]
  wire [7:0] _T_27852; // @[Mux.scala 31:69:@10507.4]
  wire [7:0] _T_27853; // @[Mux.scala 31:69:@10508.4]
  wire [7:0] _T_27854; // @[Mux.scala 31:69:@10509.4]
  wire [7:0] _T_27855; // @[Mux.scala 31:69:@10510.4]
  wire  _T_27856; // @[OneHot.scala 66:30:@10511.4]
  wire  _T_27857; // @[OneHot.scala 66:30:@10512.4]
  wire  _T_27858; // @[OneHot.scala 66:30:@10513.4]
  wire  _T_27859; // @[OneHot.scala 66:30:@10514.4]
  wire  _T_27860; // @[OneHot.scala 66:30:@10515.4]
  wire  _T_27861; // @[OneHot.scala 66:30:@10516.4]
  wire  _T_27862; // @[OneHot.scala 66:30:@10517.4]
  wire  _T_27863; // @[OneHot.scala 66:30:@10518.4]
  wire [7:0] _T_27888; // @[Mux.scala 31:69:@10528.4]
  wire [7:0] _T_27889; // @[Mux.scala 31:69:@10529.4]
  wire [7:0] _T_27890; // @[Mux.scala 31:69:@10530.4]
  wire [7:0] _T_27891; // @[Mux.scala 31:69:@10531.4]
  wire [7:0] _T_27892; // @[Mux.scala 31:69:@10532.4]
  wire [7:0] _T_27893; // @[Mux.scala 31:69:@10533.4]
  wire [7:0] _T_27894; // @[Mux.scala 31:69:@10534.4]
  wire [7:0] _T_27895; // @[Mux.scala 31:69:@10535.4]
  wire  _T_27896; // @[OneHot.scala 66:30:@10536.4]
  wire  _T_27897; // @[OneHot.scala 66:30:@10537.4]
  wire  _T_27898; // @[OneHot.scala 66:30:@10538.4]
  wire  _T_27899; // @[OneHot.scala 66:30:@10539.4]
  wire  _T_27900; // @[OneHot.scala 66:30:@10540.4]
  wire  _T_27901; // @[OneHot.scala 66:30:@10541.4]
  wire  _T_27902; // @[OneHot.scala 66:30:@10542.4]
  wire  _T_27903; // @[OneHot.scala 66:30:@10543.4]
  wire [7:0] _T_27928; // @[Mux.scala 31:69:@10553.4]
  wire [7:0] _T_27929; // @[Mux.scala 31:69:@10554.4]
  wire [7:0] _T_27930; // @[Mux.scala 31:69:@10555.4]
  wire [7:0] _T_27931; // @[Mux.scala 31:69:@10556.4]
  wire [7:0] _T_27932; // @[Mux.scala 31:69:@10557.4]
  wire [7:0] _T_27933; // @[Mux.scala 31:69:@10558.4]
  wire [7:0] _T_27934; // @[Mux.scala 31:69:@10559.4]
  wire [7:0] _T_27935; // @[Mux.scala 31:69:@10560.4]
  wire  _T_27936; // @[OneHot.scala 66:30:@10561.4]
  wire  _T_27937; // @[OneHot.scala 66:30:@10562.4]
  wire  _T_27938; // @[OneHot.scala 66:30:@10563.4]
  wire  _T_27939; // @[OneHot.scala 66:30:@10564.4]
  wire  _T_27940; // @[OneHot.scala 66:30:@10565.4]
  wire  _T_27941; // @[OneHot.scala 66:30:@10566.4]
  wire  _T_27942; // @[OneHot.scala 66:30:@10567.4]
  wire  _T_27943; // @[OneHot.scala 66:30:@10568.4]
  wire [7:0] _T_27968; // @[Mux.scala 31:69:@10578.4]
  wire [7:0] _T_27969; // @[Mux.scala 31:69:@10579.4]
  wire [7:0] _T_27970; // @[Mux.scala 31:69:@10580.4]
  wire [7:0] _T_27971; // @[Mux.scala 31:69:@10581.4]
  wire [7:0] _T_27972; // @[Mux.scala 31:69:@10582.4]
  wire [7:0] _T_27973; // @[Mux.scala 31:69:@10583.4]
  wire [7:0] _T_27974; // @[Mux.scala 31:69:@10584.4]
  wire [7:0] _T_27975; // @[Mux.scala 31:69:@10585.4]
  wire  _T_27976; // @[OneHot.scala 66:30:@10586.4]
  wire  _T_27977; // @[OneHot.scala 66:30:@10587.4]
  wire  _T_27978; // @[OneHot.scala 66:30:@10588.4]
  wire  _T_27979; // @[OneHot.scala 66:30:@10589.4]
  wire  _T_27980; // @[OneHot.scala 66:30:@10590.4]
  wire  _T_27981; // @[OneHot.scala 66:30:@10591.4]
  wire  _T_27982; // @[OneHot.scala 66:30:@10592.4]
  wire  _T_27983; // @[OneHot.scala 66:30:@10593.4]
  wire [7:0] _T_28008; // @[Mux.scala 31:69:@10603.4]
  wire [7:0] _T_28009; // @[Mux.scala 31:69:@10604.4]
  wire [7:0] _T_28010; // @[Mux.scala 31:69:@10605.4]
  wire [7:0] _T_28011; // @[Mux.scala 31:69:@10606.4]
  wire [7:0] _T_28012; // @[Mux.scala 31:69:@10607.4]
  wire [7:0] _T_28013; // @[Mux.scala 31:69:@10608.4]
  wire [7:0] _T_28014; // @[Mux.scala 31:69:@10609.4]
  wire [7:0] _T_28015; // @[Mux.scala 31:69:@10610.4]
  wire  _T_28016; // @[OneHot.scala 66:30:@10611.4]
  wire  _T_28017; // @[OneHot.scala 66:30:@10612.4]
  wire  _T_28018; // @[OneHot.scala 66:30:@10613.4]
  wire  _T_28019; // @[OneHot.scala 66:30:@10614.4]
  wire  _T_28020; // @[OneHot.scala 66:30:@10615.4]
  wire  _T_28021; // @[OneHot.scala 66:30:@10616.4]
  wire  _T_28022; // @[OneHot.scala 66:30:@10617.4]
  wire  _T_28023; // @[OneHot.scala 66:30:@10618.4]
  wire [7:0] _T_28048; // @[Mux.scala 31:69:@10628.4]
  wire [7:0] _T_28049; // @[Mux.scala 31:69:@10629.4]
  wire [7:0] _T_28050; // @[Mux.scala 31:69:@10630.4]
  wire [7:0] _T_28051; // @[Mux.scala 31:69:@10631.4]
  wire [7:0] _T_28052; // @[Mux.scala 31:69:@10632.4]
  wire [7:0] _T_28053; // @[Mux.scala 31:69:@10633.4]
  wire [7:0] _T_28054; // @[Mux.scala 31:69:@10634.4]
  wire [7:0] _T_28055; // @[Mux.scala 31:69:@10635.4]
  wire  _T_28056; // @[OneHot.scala 66:30:@10636.4]
  wire  _T_28057; // @[OneHot.scala 66:30:@10637.4]
  wire  _T_28058; // @[OneHot.scala 66:30:@10638.4]
  wire  _T_28059; // @[OneHot.scala 66:30:@10639.4]
  wire  _T_28060; // @[OneHot.scala 66:30:@10640.4]
  wire  _T_28061; // @[OneHot.scala 66:30:@10641.4]
  wire  _T_28062; // @[OneHot.scala 66:30:@10642.4]
  wire  _T_28063; // @[OneHot.scala 66:30:@10643.4]
  wire [7:0] _T_28104; // @[Mux.scala 19:72:@10659.4]
  wire [7:0] _T_28106; // @[Mux.scala 19:72:@10660.4]
  wire [7:0] _T_28113; // @[Mux.scala 19:72:@10667.4]
  wire [7:0] _T_28115; // @[Mux.scala 19:72:@10668.4]
  wire [7:0] _T_28122; // @[Mux.scala 19:72:@10675.4]
  wire [7:0] _T_28124; // @[Mux.scala 19:72:@10676.4]
  wire [7:0] _T_28131; // @[Mux.scala 19:72:@10683.4]
  wire [7:0] _T_28133; // @[Mux.scala 19:72:@10684.4]
  wire [7:0] _T_28140; // @[Mux.scala 19:72:@10691.4]
  wire [7:0] _T_28142; // @[Mux.scala 19:72:@10692.4]
  wire [7:0] _T_28149; // @[Mux.scala 19:72:@10699.4]
  wire [7:0] _T_28151; // @[Mux.scala 19:72:@10700.4]
  wire [7:0] _T_28158; // @[Mux.scala 19:72:@10707.4]
  wire [7:0] _T_28160; // @[Mux.scala 19:72:@10708.4]
  wire [7:0] _T_28167; // @[Mux.scala 19:72:@10715.4]
  wire [7:0] _T_28169; // @[Mux.scala 19:72:@10716.4]
  wire [7:0] _T_28170; // @[Mux.scala 19:72:@10717.4]
  wire [7:0] _T_28171; // @[Mux.scala 19:72:@10718.4]
  wire [7:0] _T_28172; // @[Mux.scala 19:72:@10719.4]
  wire [7:0] _T_28173; // @[Mux.scala 19:72:@10720.4]
  wire [7:0] _T_28174; // @[Mux.scala 19:72:@10721.4]
  wire [7:0] _T_28175; // @[Mux.scala 19:72:@10722.4]
  wire [7:0] _T_28176; // @[Mux.scala 19:72:@10723.4]
  wire  outputPriorityPorts_1_0; // @[Mux.scala 19:72:@10727.4]
  wire  outputPriorityPorts_1_1; // @[Mux.scala 19:72:@10729.4]
  wire  outputPriorityPorts_1_2; // @[Mux.scala 19:72:@10731.4]
  wire  outputPriorityPorts_1_3; // @[Mux.scala 19:72:@10733.4]
  wire  outputPriorityPorts_1_4; // @[Mux.scala 19:72:@10735.4]
  wire  outputPriorityPorts_1_5; // @[Mux.scala 19:72:@10737.4]
  wire  outputPriorityPorts_1_6; // @[Mux.scala 19:72:@10739.4]
  wire  outputPriorityPorts_1_7; // @[Mux.scala 19:72:@10741.4]
  wire  _T_28256; // @[LoadQueue.scala 298:83:@10752.4]
  wire  _T_28259; // @[LoadQueue.scala 298:83:@10754.4]
  wire  _T_28262; // @[LoadQueue.scala 298:83:@10756.4]
  wire  _T_28265; // @[LoadQueue.scala 298:83:@10758.4]
  wire  _T_28268; // @[LoadQueue.scala 298:83:@10760.4]
  wire  _T_28271; // @[LoadQueue.scala 298:83:@10762.4]
  wire  _T_28274; // @[LoadQueue.scala 298:83:@10764.4]
  wire  _T_28277; // @[LoadQueue.scala 298:83:@10766.4]
  wire [7:0] _T_28328; // @[Mux.scala 31:69:@10796.4]
  wire [7:0] _T_28329; // @[Mux.scala 31:69:@10797.4]
  wire [7:0] _T_28330; // @[Mux.scala 31:69:@10798.4]
  wire [7:0] _T_28331; // @[Mux.scala 31:69:@10799.4]
  wire [7:0] _T_28332; // @[Mux.scala 31:69:@10800.4]
  wire [7:0] _T_28333; // @[Mux.scala 31:69:@10801.4]
  wire [7:0] _T_28334; // @[Mux.scala 31:69:@10802.4]
  wire [7:0] _T_28335; // @[Mux.scala 31:69:@10803.4]
  wire  _T_28336; // @[OneHot.scala 66:30:@10804.4]
  wire  _T_28337; // @[OneHot.scala 66:30:@10805.4]
  wire  _T_28338; // @[OneHot.scala 66:30:@10806.4]
  wire  _T_28339; // @[OneHot.scala 66:30:@10807.4]
  wire  _T_28340; // @[OneHot.scala 66:30:@10808.4]
  wire  _T_28341; // @[OneHot.scala 66:30:@10809.4]
  wire  _T_28342; // @[OneHot.scala 66:30:@10810.4]
  wire  _T_28343; // @[OneHot.scala 66:30:@10811.4]
  wire [7:0] _T_28368; // @[Mux.scala 31:69:@10821.4]
  wire [7:0] _T_28369; // @[Mux.scala 31:69:@10822.4]
  wire [7:0] _T_28370; // @[Mux.scala 31:69:@10823.4]
  wire [7:0] _T_28371; // @[Mux.scala 31:69:@10824.4]
  wire [7:0] _T_28372; // @[Mux.scala 31:69:@10825.4]
  wire [7:0] _T_28373; // @[Mux.scala 31:69:@10826.4]
  wire [7:0] _T_28374; // @[Mux.scala 31:69:@10827.4]
  wire [7:0] _T_28375; // @[Mux.scala 31:69:@10828.4]
  wire  _T_28376; // @[OneHot.scala 66:30:@10829.4]
  wire  _T_28377; // @[OneHot.scala 66:30:@10830.4]
  wire  _T_28378; // @[OneHot.scala 66:30:@10831.4]
  wire  _T_28379; // @[OneHot.scala 66:30:@10832.4]
  wire  _T_28380; // @[OneHot.scala 66:30:@10833.4]
  wire  _T_28381; // @[OneHot.scala 66:30:@10834.4]
  wire  _T_28382; // @[OneHot.scala 66:30:@10835.4]
  wire  _T_28383; // @[OneHot.scala 66:30:@10836.4]
  wire [7:0] _T_28408; // @[Mux.scala 31:69:@10846.4]
  wire [7:0] _T_28409; // @[Mux.scala 31:69:@10847.4]
  wire [7:0] _T_28410; // @[Mux.scala 31:69:@10848.4]
  wire [7:0] _T_28411; // @[Mux.scala 31:69:@10849.4]
  wire [7:0] _T_28412; // @[Mux.scala 31:69:@10850.4]
  wire [7:0] _T_28413; // @[Mux.scala 31:69:@10851.4]
  wire [7:0] _T_28414; // @[Mux.scala 31:69:@10852.4]
  wire [7:0] _T_28415; // @[Mux.scala 31:69:@10853.4]
  wire  _T_28416; // @[OneHot.scala 66:30:@10854.4]
  wire  _T_28417; // @[OneHot.scala 66:30:@10855.4]
  wire  _T_28418; // @[OneHot.scala 66:30:@10856.4]
  wire  _T_28419; // @[OneHot.scala 66:30:@10857.4]
  wire  _T_28420; // @[OneHot.scala 66:30:@10858.4]
  wire  _T_28421; // @[OneHot.scala 66:30:@10859.4]
  wire  _T_28422; // @[OneHot.scala 66:30:@10860.4]
  wire  _T_28423; // @[OneHot.scala 66:30:@10861.4]
  wire [7:0] _T_28448; // @[Mux.scala 31:69:@10871.4]
  wire [7:0] _T_28449; // @[Mux.scala 31:69:@10872.4]
  wire [7:0] _T_28450; // @[Mux.scala 31:69:@10873.4]
  wire [7:0] _T_28451; // @[Mux.scala 31:69:@10874.4]
  wire [7:0] _T_28452; // @[Mux.scala 31:69:@10875.4]
  wire [7:0] _T_28453; // @[Mux.scala 31:69:@10876.4]
  wire [7:0] _T_28454; // @[Mux.scala 31:69:@10877.4]
  wire [7:0] _T_28455; // @[Mux.scala 31:69:@10878.4]
  wire  _T_28456; // @[OneHot.scala 66:30:@10879.4]
  wire  _T_28457; // @[OneHot.scala 66:30:@10880.4]
  wire  _T_28458; // @[OneHot.scala 66:30:@10881.4]
  wire  _T_28459; // @[OneHot.scala 66:30:@10882.4]
  wire  _T_28460; // @[OneHot.scala 66:30:@10883.4]
  wire  _T_28461; // @[OneHot.scala 66:30:@10884.4]
  wire  _T_28462; // @[OneHot.scala 66:30:@10885.4]
  wire  _T_28463; // @[OneHot.scala 66:30:@10886.4]
  wire [7:0] _T_28488; // @[Mux.scala 31:69:@10896.4]
  wire [7:0] _T_28489; // @[Mux.scala 31:69:@10897.4]
  wire [7:0] _T_28490; // @[Mux.scala 31:69:@10898.4]
  wire [7:0] _T_28491; // @[Mux.scala 31:69:@10899.4]
  wire [7:0] _T_28492; // @[Mux.scala 31:69:@10900.4]
  wire [7:0] _T_28493; // @[Mux.scala 31:69:@10901.4]
  wire [7:0] _T_28494; // @[Mux.scala 31:69:@10902.4]
  wire [7:0] _T_28495; // @[Mux.scala 31:69:@10903.4]
  wire  _T_28496; // @[OneHot.scala 66:30:@10904.4]
  wire  _T_28497; // @[OneHot.scala 66:30:@10905.4]
  wire  _T_28498; // @[OneHot.scala 66:30:@10906.4]
  wire  _T_28499; // @[OneHot.scala 66:30:@10907.4]
  wire  _T_28500; // @[OneHot.scala 66:30:@10908.4]
  wire  _T_28501; // @[OneHot.scala 66:30:@10909.4]
  wire  _T_28502; // @[OneHot.scala 66:30:@10910.4]
  wire  _T_28503; // @[OneHot.scala 66:30:@10911.4]
  wire [7:0] _T_28528; // @[Mux.scala 31:69:@10921.4]
  wire [7:0] _T_28529; // @[Mux.scala 31:69:@10922.4]
  wire [7:0] _T_28530; // @[Mux.scala 31:69:@10923.4]
  wire [7:0] _T_28531; // @[Mux.scala 31:69:@10924.4]
  wire [7:0] _T_28532; // @[Mux.scala 31:69:@10925.4]
  wire [7:0] _T_28533; // @[Mux.scala 31:69:@10926.4]
  wire [7:0] _T_28534; // @[Mux.scala 31:69:@10927.4]
  wire [7:0] _T_28535; // @[Mux.scala 31:69:@10928.4]
  wire  _T_28536; // @[OneHot.scala 66:30:@10929.4]
  wire  _T_28537; // @[OneHot.scala 66:30:@10930.4]
  wire  _T_28538; // @[OneHot.scala 66:30:@10931.4]
  wire  _T_28539; // @[OneHot.scala 66:30:@10932.4]
  wire  _T_28540; // @[OneHot.scala 66:30:@10933.4]
  wire  _T_28541; // @[OneHot.scala 66:30:@10934.4]
  wire  _T_28542; // @[OneHot.scala 66:30:@10935.4]
  wire  _T_28543; // @[OneHot.scala 66:30:@10936.4]
  wire [7:0] _T_28568; // @[Mux.scala 31:69:@10946.4]
  wire [7:0] _T_28569; // @[Mux.scala 31:69:@10947.4]
  wire [7:0] _T_28570; // @[Mux.scala 31:69:@10948.4]
  wire [7:0] _T_28571; // @[Mux.scala 31:69:@10949.4]
  wire [7:0] _T_28572; // @[Mux.scala 31:69:@10950.4]
  wire [7:0] _T_28573; // @[Mux.scala 31:69:@10951.4]
  wire [7:0] _T_28574; // @[Mux.scala 31:69:@10952.4]
  wire [7:0] _T_28575; // @[Mux.scala 31:69:@10953.4]
  wire  _T_28576; // @[OneHot.scala 66:30:@10954.4]
  wire  _T_28577; // @[OneHot.scala 66:30:@10955.4]
  wire  _T_28578; // @[OneHot.scala 66:30:@10956.4]
  wire  _T_28579; // @[OneHot.scala 66:30:@10957.4]
  wire  _T_28580; // @[OneHot.scala 66:30:@10958.4]
  wire  _T_28581; // @[OneHot.scala 66:30:@10959.4]
  wire  _T_28582; // @[OneHot.scala 66:30:@10960.4]
  wire  _T_28583; // @[OneHot.scala 66:30:@10961.4]
  wire [7:0] _T_28608; // @[Mux.scala 31:69:@10971.4]
  wire [7:0] _T_28609; // @[Mux.scala 31:69:@10972.4]
  wire [7:0] _T_28610; // @[Mux.scala 31:69:@10973.4]
  wire [7:0] _T_28611; // @[Mux.scala 31:69:@10974.4]
  wire [7:0] _T_28612; // @[Mux.scala 31:69:@10975.4]
  wire [7:0] _T_28613; // @[Mux.scala 31:69:@10976.4]
  wire [7:0] _T_28614; // @[Mux.scala 31:69:@10977.4]
  wire [7:0] _T_28615; // @[Mux.scala 31:69:@10978.4]
  wire  _T_28616; // @[OneHot.scala 66:30:@10979.4]
  wire  _T_28617; // @[OneHot.scala 66:30:@10980.4]
  wire  _T_28618; // @[OneHot.scala 66:30:@10981.4]
  wire  _T_28619; // @[OneHot.scala 66:30:@10982.4]
  wire  _T_28620; // @[OneHot.scala 66:30:@10983.4]
  wire  _T_28621; // @[OneHot.scala 66:30:@10984.4]
  wire  _T_28622; // @[OneHot.scala 66:30:@10985.4]
  wire  _T_28623; // @[OneHot.scala 66:30:@10986.4]
  wire [7:0] _T_28664; // @[Mux.scala 19:72:@11002.4]
  wire [7:0] _T_28666; // @[Mux.scala 19:72:@11003.4]
  wire [7:0] _T_28673; // @[Mux.scala 19:72:@11010.4]
  wire [7:0] _T_28675; // @[Mux.scala 19:72:@11011.4]
  wire [7:0] _T_28682; // @[Mux.scala 19:72:@11018.4]
  wire [7:0] _T_28684; // @[Mux.scala 19:72:@11019.4]
  wire [7:0] _T_28691; // @[Mux.scala 19:72:@11026.4]
  wire [7:0] _T_28693; // @[Mux.scala 19:72:@11027.4]
  wire [7:0] _T_28700; // @[Mux.scala 19:72:@11034.4]
  wire [7:0] _T_28702; // @[Mux.scala 19:72:@11035.4]
  wire [7:0] _T_28709; // @[Mux.scala 19:72:@11042.4]
  wire [7:0] _T_28711; // @[Mux.scala 19:72:@11043.4]
  wire [7:0] _T_28718; // @[Mux.scala 19:72:@11050.4]
  wire [7:0] _T_28720; // @[Mux.scala 19:72:@11051.4]
  wire [7:0] _T_28727; // @[Mux.scala 19:72:@11058.4]
  wire [7:0] _T_28729; // @[Mux.scala 19:72:@11059.4]
  wire [7:0] _T_28730; // @[Mux.scala 19:72:@11060.4]
  wire [7:0] _T_28731; // @[Mux.scala 19:72:@11061.4]
  wire [7:0] _T_28732; // @[Mux.scala 19:72:@11062.4]
  wire [7:0] _T_28733; // @[Mux.scala 19:72:@11063.4]
  wire [7:0] _T_28734; // @[Mux.scala 19:72:@11064.4]
  wire [7:0] _T_28735; // @[Mux.scala 19:72:@11065.4]
  wire [7:0] _T_28736; // @[Mux.scala 19:72:@11066.4]
  wire  inputPriorityPorts_2_0; // @[Mux.scala 19:72:@11070.4]
  wire  inputPriorityPorts_2_1; // @[Mux.scala 19:72:@11072.4]
  wire  inputPriorityPorts_2_2; // @[Mux.scala 19:72:@11074.4]
  wire  inputPriorityPorts_2_3; // @[Mux.scala 19:72:@11076.4]
  wire  inputPriorityPorts_2_4; // @[Mux.scala 19:72:@11078.4]
  wire  inputPriorityPorts_2_5; // @[Mux.scala 19:72:@11080.4]
  wire  inputPriorityPorts_2_6; // @[Mux.scala 19:72:@11082.4]
  wire  inputPriorityPorts_2_7; // @[Mux.scala 19:72:@11084.4]
  wire [7:0] _T_28850; // @[Mux.scala 31:69:@11114.4]
  wire [7:0] _T_28851; // @[Mux.scala 31:69:@11115.4]
  wire [7:0] _T_28852; // @[Mux.scala 31:69:@11116.4]
  wire [7:0] _T_28853; // @[Mux.scala 31:69:@11117.4]
  wire [7:0] _T_28854; // @[Mux.scala 31:69:@11118.4]
  wire [7:0] _T_28855; // @[Mux.scala 31:69:@11119.4]
  wire [7:0] _T_28856; // @[Mux.scala 31:69:@11120.4]
  wire [7:0] _T_28857; // @[Mux.scala 31:69:@11121.4]
  wire  _T_28858; // @[OneHot.scala 66:30:@11122.4]
  wire  _T_28859; // @[OneHot.scala 66:30:@11123.4]
  wire  _T_28860; // @[OneHot.scala 66:30:@11124.4]
  wire  _T_28861; // @[OneHot.scala 66:30:@11125.4]
  wire  _T_28862; // @[OneHot.scala 66:30:@11126.4]
  wire  _T_28863; // @[OneHot.scala 66:30:@11127.4]
  wire  _T_28864; // @[OneHot.scala 66:30:@11128.4]
  wire  _T_28865; // @[OneHot.scala 66:30:@11129.4]
  wire [7:0] _T_28890; // @[Mux.scala 31:69:@11139.4]
  wire [7:0] _T_28891; // @[Mux.scala 31:69:@11140.4]
  wire [7:0] _T_28892; // @[Mux.scala 31:69:@11141.4]
  wire [7:0] _T_28893; // @[Mux.scala 31:69:@11142.4]
  wire [7:0] _T_28894; // @[Mux.scala 31:69:@11143.4]
  wire [7:0] _T_28895; // @[Mux.scala 31:69:@11144.4]
  wire [7:0] _T_28896; // @[Mux.scala 31:69:@11145.4]
  wire [7:0] _T_28897; // @[Mux.scala 31:69:@11146.4]
  wire  _T_28898; // @[OneHot.scala 66:30:@11147.4]
  wire  _T_28899; // @[OneHot.scala 66:30:@11148.4]
  wire  _T_28900; // @[OneHot.scala 66:30:@11149.4]
  wire  _T_28901; // @[OneHot.scala 66:30:@11150.4]
  wire  _T_28902; // @[OneHot.scala 66:30:@11151.4]
  wire  _T_28903; // @[OneHot.scala 66:30:@11152.4]
  wire  _T_28904; // @[OneHot.scala 66:30:@11153.4]
  wire  _T_28905; // @[OneHot.scala 66:30:@11154.4]
  wire [7:0] _T_28930; // @[Mux.scala 31:69:@11164.4]
  wire [7:0] _T_28931; // @[Mux.scala 31:69:@11165.4]
  wire [7:0] _T_28932; // @[Mux.scala 31:69:@11166.4]
  wire [7:0] _T_28933; // @[Mux.scala 31:69:@11167.4]
  wire [7:0] _T_28934; // @[Mux.scala 31:69:@11168.4]
  wire [7:0] _T_28935; // @[Mux.scala 31:69:@11169.4]
  wire [7:0] _T_28936; // @[Mux.scala 31:69:@11170.4]
  wire [7:0] _T_28937; // @[Mux.scala 31:69:@11171.4]
  wire  _T_28938; // @[OneHot.scala 66:30:@11172.4]
  wire  _T_28939; // @[OneHot.scala 66:30:@11173.4]
  wire  _T_28940; // @[OneHot.scala 66:30:@11174.4]
  wire  _T_28941; // @[OneHot.scala 66:30:@11175.4]
  wire  _T_28942; // @[OneHot.scala 66:30:@11176.4]
  wire  _T_28943; // @[OneHot.scala 66:30:@11177.4]
  wire  _T_28944; // @[OneHot.scala 66:30:@11178.4]
  wire  _T_28945; // @[OneHot.scala 66:30:@11179.4]
  wire [7:0] _T_28970; // @[Mux.scala 31:69:@11189.4]
  wire [7:0] _T_28971; // @[Mux.scala 31:69:@11190.4]
  wire [7:0] _T_28972; // @[Mux.scala 31:69:@11191.4]
  wire [7:0] _T_28973; // @[Mux.scala 31:69:@11192.4]
  wire [7:0] _T_28974; // @[Mux.scala 31:69:@11193.4]
  wire [7:0] _T_28975; // @[Mux.scala 31:69:@11194.4]
  wire [7:0] _T_28976; // @[Mux.scala 31:69:@11195.4]
  wire [7:0] _T_28977; // @[Mux.scala 31:69:@11196.4]
  wire  _T_28978; // @[OneHot.scala 66:30:@11197.4]
  wire  _T_28979; // @[OneHot.scala 66:30:@11198.4]
  wire  _T_28980; // @[OneHot.scala 66:30:@11199.4]
  wire  _T_28981; // @[OneHot.scala 66:30:@11200.4]
  wire  _T_28982; // @[OneHot.scala 66:30:@11201.4]
  wire  _T_28983; // @[OneHot.scala 66:30:@11202.4]
  wire  _T_28984; // @[OneHot.scala 66:30:@11203.4]
  wire  _T_28985; // @[OneHot.scala 66:30:@11204.4]
  wire [7:0] _T_29010; // @[Mux.scala 31:69:@11214.4]
  wire [7:0] _T_29011; // @[Mux.scala 31:69:@11215.4]
  wire [7:0] _T_29012; // @[Mux.scala 31:69:@11216.4]
  wire [7:0] _T_29013; // @[Mux.scala 31:69:@11217.4]
  wire [7:0] _T_29014; // @[Mux.scala 31:69:@11218.4]
  wire [7:0] _T_29015; // @[Mux.scala 31:69:@11219.4]
  wire [7:0] _T_29016; // @[Mux.scala 31:69:@11220.4]
  wire [7:0] _T_29017; // @[Mux.scala 31:69:@11221.4]
  wire  _T_29018; // @[OneHot.scala 66:30:@11222.4]
  wire  _T_29019; // @[OneHot.scala 66:30:@11223.4]
  wire  _T_29020; // @[OneHot.scala 66:30:@11224.4]
  wire  _T_29021; // @[OneHot.scala 66:30:@11225.4]
  wire  _T_29022; // @[OneHot.scala 66:30:@11226.4]
  wire  _T_29023; // @[OneHot.scala 66:30:@11227.4]
  wire  _T_29024; // @[OneHot.scala 66:30:@11228.4]
  wire  _T_29025; // @[OneHot.scala 66:30:@11229.4]
  wire [7:0] _T_29050; // @[Mux.scala 31:69:@11239.4]
  wire [7:0] _T_29051; // @[Mux.scala 31:69:@11240.4]
  wire [7:0] _T_29052; // @[Mux.scala 31:69:@11241.4]
  wire [7:0] _T_29053; // @[Mux.scala 31:69:@11242.4]
  wire [7:0] _T_29054; // @[Mux.scala 31:69:@11243.4]
  wire [7:0] _T_29055; // @[Mux.scala 31:69:@11244.4]
  wire [7:0] _T_29056; // @[Mux.scala 31:69:@11245.4]
  wire [7:0] _T_29057; // @[Mux.scala 31:69:@11246.4]
  wire  _T_29058; // @[OneHot.scala 66:30:@11247.4]
  wire  _T_29059; // @[OneHot.scala 66:30:@11248.4]
  wire  _T_29060; // @[OneHot.scala 66:30:@11249.4]
  wire  _T_29061; // @[OneHot.scala 66:30:@11250.4]
  wire  _T_29062; // @[OneHot.scala 66:30:@11251.4]
  wire  _T_29063; // @[OneHot.scala 66:30:@11252.4]
  wire  _T_29064; // @[OneHot.scala 66:30:@11253.4]
  wire  _T_29065; // @[OneHot.scala 66:30:@11254.4]
  wire [7:0] _T_29090; // @[Mux.scala 31:69:@11264.4]
  wire [7:0] _T_29091; // @[Mux.scala 31:69:@11265.4]
  wire [7:0] _T_29092; // @[Mux.scala 31:69:@11266.4]
  wire [7:0] _T_29093; // @[Mux.scala 31:69:@11267.4]
  wire [7:0] _T_29094; // @[Mux.scala 31:69:@11268.4]
  wire [7:0] _T_29095; // @[Mux.scala 31:69:@11269.4]
  wire [7:0] _T_29096; // @[Mux.scala 31:69:@11270.4]
  wire [7:0] _T_29097; // @[Mux.scala 31:69:@11271.4]
  wire  _T_29098; // @[OneHot.scala 66:30:@11272.4]
  wire  _T_29099; // @[OneHot.scala 66:30:@11273.4]
  wire  _T_29100; // @[OneHot.scala 66:30:@11274.4]
  wire  _T_29101; // @[OneHot.scala 66:30:@11275.4]
  wire  _T_29102; // @[OneHot.scala 66:30:@11276.4]
  wire  _T_29103; // @[OneHot.scala 66:30:@11277.4]
  wire  _T_29104; // @[OneHot.scala 66:30:@11278.4]
  wire  _T_29105; // @[OneHot.scala 66:30:@11279.4]
  wire [7:0] _T_29130; // @[Mux.scala 31:69:@11289.4]
  wire [7:0] _T_29131; // @[Mux.scala 31:69:@11290.4]
  wire [7:0] _T_29132; // @[Mux.scala 31:69:@11291.4]
  wire [7:0] _T_29133; // @[Mux.scala 31:69:@11292.4]
  wire [7:0] _T_29134; // @[Mux.scala 31:69:@11293.4]
  wire [7:0] _T_29135; // @[Mux.scala 31:69:@11294.4]
  wire [7:0] _T_29136; // @[Mux.scala 31:69:@11295.4]
  wire [7:0] _T_29137; // @[Mux.scala 31:69:@11296.4]
  wire  _T_29138; // @[OneHot.scala 66:30:@11297.4]
  wire  _T_29139; // @[OneHot.scala 66:30:@11298.4]
  wire  _T_29140; // @[OneHot.scala 66:30:@11299.4]
  wire  _T_29141; // @[OneHot.scala 66:30:@11300.4]
  wire  _T_29142; // @[OneHot.scala 66:30:@11301.4]
  wire  _T_29143; // @[OneHot.scala 66:30:@11302.4]
  wire  _T_29144; // @[OneHot.scala 66:30:@11303.4]
  wire  _T_29145; // @[OneHot.scala 66:30:@11304.4]
  wire [7:0] _T_29186; // @[Mux.scala 19:72:@11320.4]
  wire [7:0] _T_29188; // @[Mux.scala 19:72:@11321.4]
  wire [7:0] _T_29195; // @[Mux.scala 19:72:@11328.4]
  wire [7:0] _T_29197; // @[Mux.scala 19:72:@11329.4]
  wire [7:0] _T_29204; // @[Mux.scala 19:72:@11336.4]
  wire [7:0] _T_29206; // @[Mux.scala 19:72:@11337.4]
  wire [7:0] _T_29213; // @[Mux.scala 19:72:@11344.4]
  wire [7:0] _T_29215; // @[Mux.scala 19:72:@11345.4]
  wire [7:0] _T_29222; // @[Mux.scala 19:72:@11352.4]
  wire [7:0] _T_29224; // @[Mux.scala 19:72:@11353.4]
  wire [7:0] _T_29231; // @[Mux.scala 19:72:@11360.4]
  wire [7:0] _T_29233; // @[Mux.scala 19:72:@11361.4]
  wire [7:0] _T_29240; // @[Mux.scala 19:72:@11368.4]
  wire [7:0] _T_29242; // @[Mux.scala 19:72:@11369.4]
  wire [7:0] _T_29249; // @[Mux.scala 19:72:@11376.4]
  wire [7:0] _T_29251; // @[Mux.scala 19:72:@11377.4]
  wire [7:0] _T_29252; // @[Mux.scala 19:72:@11378.4]
  wire [7:0] _T_29253; // @[Mux.scala 19:72:@11379.4]
  wire [7:0] _T_29254; // @[Mux.scala 19:72:@11380.4]
  wire [7:0] _T_29255; // @[Mux.scala 19:72:@11381.4]
  wire [7:0] _T_29256; // @[Mux.scala 19:72:@11382.4]
  wire [7:0] _T_29257; // @[Mux.scala 19:72:@11383.4]
  wire [7:0] _T_29258; // @[Mux.scala 19:72:@11384.4]
  wire  outputPriorityPorts_2_0; // @[Mux.scala 19:72:@11388.4]
  wire  outputPriorityPorts_2_1; // @[Mux.scala 19:72:@11390.4]
  wire  outputPriorityPorts_2_2; // @[Mux.scala 19:72:@11392.4]
  wire  outputPriorityPorts_2_3; // @[Mux.scala 19:72:@11394.4]
  wire  outputPriorityPorts_2_4; // @[Mux.scala 19:72:@11396.4]
  wire  outputPriorityPorts_2_5; // @[Mux.scala 19:72:@11398.4]
  wire  outputPriorityPorts_2_6; // @[Mux.scala 19:72:@11400.4]
  wire  outputPriorityPorts_2_7; // @[Mux.scala 19:72:@11402.4]
  wire  _T_29338; // @[LoadQueue.scala 298:83:@11413.4]
  wire  _T_29341; // @[LoadQueue.scala 298:83:@11415.4]
  wire  _T_29344; // @[LoadQueue.scala 298:83:@11417.4]
  wire  _T_29347; // @[LoadQueue.scala 298:83:@11419.4]
  wire  _T_29350; // @[LoadQueue.scala 298:83:@11421.4]
  wire  _T_29353; // @[LoadQueue.scala 298:83:@11423.4]
  wire  _T_29356; // @[LoadQueue.scala 298:83:@11425.4]
  wire  _T_29359; // @[LoadQueue.scala 298:83:@11427.4]
  wire [7:0] _T_29410; // @[Mux.scala 31:69:@11457.4]
  wire [7:0] _T_29411; // @[Mux.scala 31:69:@11458.4]
  wire [7:0] _T_29412; // @[Mux.scala 31:69:@11459.4]
  wire [7:0] _T_29413; // @[Mux.scala 31:69:@11460.4]
  wire [7:0] _T_29414; // @[Mux.scala 31:69:@11461.4]
  wire [7:0] _T_29415; // @[Mux.scala 31:69:@11462.4]
  wire [7:0] _T_29416; // @[Mux.scala 31:69:@11463.4]
  wire [7:0] _T_29417; // @[Mux.scala 31:69:@11464.4]
  wire  _T_29418; // @[OneHot.scala 66:30:@11465.4]
  wire  _T_29419; // @[OneHot.scala 66:30:@11466.4]
  wire  _T_29420; // @[OneHot.scala 66:30:@11467.4]
  wire  _T_29421; // @[OneHot.scala 66:30:@11468.4]
  wire  _T_29422; // @[OneHot.scala 66:30:@11469.4]
  wire  _T_29423; // @[OneHot.scala 66:30:@11470.4]
  wire  _T_29424; // @[OneHot.scala 66:30:@11471.4]
  wire  _T_29425; // @[OneHot.scala 66:30:@11472.4]
  wire [7:0] _T_29450; // @[Mux.scala 31:69:@11482.4]
  wire [7:0] _T_29451; // @[Mux.scala 31:69:@11483.4]
  wire [7:0] _T_29452; // @[Mux.scala 31:69:@11484.4]
  wire [7:0] _T_29453; // @[Mux.scala 31:69:@11485.4]
  wire [7:0] _T_29454; // @[Mux.scala 31:69:@11486.4]
  wire [7:0] _T_29455; // @[Mux.scala 31:69:@11487.4]
  wire [7:0] _T_29456; // @[Mux.scala 31:69:@11488.4]
  wire [7:0] _T_29457; // @[Mux.scala 31:69:@11489.4]
  wire  _T_29458; // @[OneHot.scala 66:30:@11490.4]
  wire  _T_29459; // @[OneHot.scala 66:30:@11491.4]
  wire  _T_29460; // @[OneHot.scala 66:30:@11492.4]
  wire  _T_29461; // @[OneHot.scala 66:30:@11493.4]
  wire  _T_29462; // @[OneHot.scala 66:30:@11494.4]
  wire  _T_29463; // @[OneHot.scala 66:30:@11495.4]
  wire  _T_29464; // @[OneHot.scala 66:30:@11496.4]
  wire  _T_29465; // @[OneHot.scala 66:30:@11497.4]
  wire [7:0] _T_29490; // @[Mux.scala 31:69:@11507.4]
  wire [7:0] _T_29491; // @[Mux.scala 31:69:@11508.4]
  wire [7:0] _T_29492; // @[Mux.scala 31:69:@11509.4]
  wire [7:0] _T_29493; // @[Mux.scala 31:69:@11510.4]
  wire [7:0] _T_29494; // @[Mux.scala 31:69:@11511.4]
  wire [7:0] _T_29495; // @[Mux.scala 31:69:@11512.4]
  wire [7:0] _T_29496; // @[Mux.scala 31:69:@11513.4]
  wire [7:0] _T_29497; // @[Mux.scala 31:69:@11514.4]
  wire  _T_29498; // @[OneHot.scala 66:30:@11515.4]
  wire  _T_29499; // @[OneHot.scala 66:30:@11516.4]
  wire  _T_29500; // @[OneHot.scala 66:30:@11517.4]
  wire  _T_29501; // @[OneHot.scala 66:30:@11518.4]
  wire  _T_29502; // @[OneHot.scala 66:30:@11519.4]
  wire  _T_29503; // @[OneHot.scala 66:30:@11520.4]
  wire  _T_29504; // @[OneHot.scala 66:30:@11521.4]
  wire  _T_29505; // @[OneHot.scala 66:30:@11522.4]
  wire [7:0] _T_29530; // @[Mux.scala 31:69:@11532.4]
  wire [7:0] _T_29531; // @[Mux.scala 31:69:@11533.4]
  wire [7:0] _T_29532; // @[Mux.scala 31:69:@11534.4]
  wire [7:0] _T_29533; // @[Mux.scala 31:69:@11535.4]
  wire [7:0] _T_29534; // @[Mux.scala 31:69:@11536.4]
  wire [7:0] _T_29535; // @[Mux.scala 31:69:@11537.4]
  wire [7:0] _T_29536; // @[Mux.scala 31:69:@11538.4]
  wire [7:0] _T_29537; // @[Mux.scala 31:69:@11539.4]
  wire  _T_29538; // @[OneHot.scala 66:30:@11540.4]
  wire  _T_29539; // @[OneHot.scala 66:30:@11541.4]
  wire  _T_29540; // @[OneHot.scala 66:30:@11542.4]
  wire  _T_29541; // @[OneHot.scala 66:30:@11543.4]
  wire  _T_29542; // @[OneHot.scala 66:30:@11544.4]
  wire  _T_29543; // @[OneHot.scala 66:30:@11545.4]
  wire  _T_29544; // @[OneHot.scala 66:30:@11546.4]
  wire  _T_29545; // @[OneHot.scala 66:30:@11547.4]
  wire [7:0] _T_29570; // @[Mux.scala 31:69:@11557.4]
  wire [7:0] _T_29571; // @[Mux.scala 31:69:@11558.4]
  wire [7:0] _T_29572; // @[Mux.scala 31:69:@11559.4]
  wire [7:0] _T_29573; // @[Mux.scala 31:69:@11560.4]
  wire [7:0] _T_29574; // @[Mux.scala 31:69:@11561.4]
  wire [7:0] _T_29575; // @[Mux.scala 31:69:@11562.4]
  wire [7:0] _T_29576; // @[Mux.scala 31:69:@11563.4]
  wire [7:0] _T_29577; // @[Mux.scala 31:69:@11564.4]
  wire  _T_29578; // @[OneHot.scala 66:30:@11565.4]
  wire  _T_29579; // @[OneHot.scala 66:30:@11566.4]
  wire  _T_29580; // @[OneHot.scala 66:30:@11567.4]
  wire  _T_29581; // @[OneHot.scala 66:30:@11568.4]
  wire  _T_29582; // @[OneHot.scala 66:30:@11569.4]
  wire  _T_29583; // @[OneHot.scala 66:30:@11570.4]
  wire  _T_29584; // @[OneHot.scala 66:30:@11571.4]
  wire  _T_29585; // @[OneHot.scala 66:30:@11572.4]
  wire [7:0] _T_29610; // @[Mux.scala 31:69:@11582.4]
  wire [7:0] _T_29611; // @[Mux.scala 31:69:@11583.4]
  wire [7:0] _T_29612; // @[Mux.scala 31:69:@11584.4]
  wire [7:0] _T_29613; // @[Mux.scala 31:69:@11585.4]
  wire [7:0] _T_29614; // @[Mux.scala 31:69:@11586.4]
  wire [7:0] _T_29615; // @[Mux.scala 31:69:@11587.4]
  wire [7:0] _T_29616; // @[Mux.scala 31:69:@11588.4]
  wire [7:0] _T_29617; // @[Mux.scala 31:69:@11589.4]
  wire  _T_29618; // @[OneHot.scala 66:30:@11590.4]
  wire  _T_29619; // @[OneHot.scala 66:30:@11591.4]
  wire  _T_29620; // @[OneHot.scala 66:30:@11592.4]
  wire  _T_29621; // @[OneHot.scala 66:30:@11593.4]
  wire  _T_29622; // @[OneHot.scala 66:30:@11594.4]
  wire  _T_29623; // @[OneHot.scala 66:30:@11595.4]
  wire  _T_29624; // @[OneHot.scala 66:30:@11596.4]
  wire  _T_29625; // @[OneHot.scala 66:30:@11597.4]
  wire [7:0] _T_29650; // @[Mux.scala 31:69:@11607.4]
  wire [7:0] _T_29651; // @[Mux.scala 31:69:@11608.4]
  wire [7:0] _T_29652; // @[Mux.scala 31:69:@11609.4]
  wire [7:0] _T_29653; // @[Mux.scala 31:69:@11610.4]
  wire [7:0] _T_29654; // @[Mux.scala 31:69:@11611.4]
  wire [7:0] _T_29655; // @[Mux.scala 31:69:@11612.4]
  wire [7:0] _T_29656; // @[Mux.scala 31:69:@11613.4]
  wire [7:0] _T_29657; // @[Mux.scala 31:69:@11614.4]
  wire  _T_29658; // @[OneHot.scala 66:30:@11615.4]
  wire  _T_29659; // @[OneHot.scala 66:30:@11616.4]
  wire  _T_29660; // @[OneHot.scala 66:30:@11617.4]
  wire  _T_29661; // @[OneHot.scala 66:30:@11618.4]
  wire  _T_29662; // @[OneHot.scala 66:30:@11619.4]
  wire  _T_29663; // @[OneHot.scala 66:30:@11620.4]
  wire  _T_29664; // @[OneHot.scala 66:30:@11621.4]
  wire  _T_29665; // @[OneHot.scala 66:30:@11622.4]
  wire [7:0] _T_29690; // @[Mux.scala 31:69:@11632.4]
  wire [7:0] _T_29691; // @[Mux.scala 31:69:@11633.4]
  wire [7:0] _T_29692; // @[Mux.scala 31:69:@11634.4]
  wire [7:0] _T_29693; // @[Mux.scala 31:69:@11635.4]
  wire [7:0] _T_29694; // @[Mux.scala 31:69:@11636.4]
  wire [7:0] _T_29695; // @[Mux.scala 31:69:@11637.4]
  wire [7:0] _T_29696; // @[Mux.scala 31:69:@11638.4]
  wire [7:0] _T_29697; // @[Mux.scala 31:69:@11639.4]
  wire  _T_29698; // @[OneHot.scala 66:30:@11640.4]
  wire  _T_29699; // @[OneHot.scala 66:30:@11641.4]
  wire  _T_29700; // @[OneHot.scala 66:30:@11642.4]
  wire  _T_29701; // @[OneHot.scala 66:30:@11643.4]
  wire  _T_29702; // @[OneHot.scala 66:30:@11644.4]
  wire  _T_29703; // @[OneHot.scala 66:30:@11645.4]
  wire  _T_29704; // @[OneHot.scala 66:30:@11646.4]
  wire  _T_29705; // @[OneHot.scala 66:30:@11647.4]
  wire [7:0] _T_29746; // @[Mux.scala 19:72:@11663.4]
  wire [7:0] _T_29748; // @[Mux.scala 19:72:@11664.4]
  wire [7:0] _T_29755; // @[Mux.scala 19:72:@11671.4]
  wire [7:0] _T_29757; // @[Mux.scala 19:72:@11672.4]
  wire [7:0] _T_29764; // @[Mux.scala 19:72:@11679.4]
  wire [7:0] _T_29766; // @[Mux.scala 19:72:@11680.4]
  wire [7:0] _T_29773; // @[Mux.scala 19:72:@11687.4]
  wire [7:0] _T_29775; // @[Mux.scala 19:72:@11688.4]
  wire [7:0] _T_29782; // @[Mux.scala 19:72:@11695.4]
  wire [7:0] _T_29784; // @[Mux.scala 19:72:@11696.4]
  wire [7:0] _T_29791; // @[Mux.scala 19:72:@11703.4]
  wire [7:0] _T_29793; // @[Mux.scala 19:72:@11704.4]
  wire [7:0] _T_29800; // @[Mux.scala 19:72:@11711.4]
  wire [7:0] _T_29802; // @[Mux.scala 19:72:@11712.4]
  wire [7:0] _T_29809; // @[Mux.scala 19:72:@11719.4]
  wire [7:0] _T_29811; // @[Mux.scala 19:72:@11720.4]
  wire [7:0] _T_29812; // @[Mux.scala 19:72:@11721.4]
  wire [7:0] _T_29813; // @[Mux.scala 19:72:@11722.4]
  wire [7:0] _T_29814; // @[Mux.scala 19:72:@11723.4]
  wire [7:0] _T_29815; // @[Mux.scala 19:72:@11724.4]
  wire [7:0] _T_29816; // @[Mux.scala 19:72:@11725.4]
  wire [7:0] _T_29817; // @[Mux.scala 19:72:@11726.4]
  wire [7:0] _T_29818; // @[Mux.scala 19:72:@11727.4]
  wire  inputPriorityPorts_3_0; // @[Mux.scala 19:72:@11731.4]
  wire  inputPriorityPorts_3_1; // @[Mux.scala 19:72:@11733.4]
  wire  inputPriorityPorts_3_2; // @[Mux.scala 19:72:@11735.4]
  wire  inputPriorityPorts_3_3; // @[Mux.scala 19:72:@11737.4]
  wire  inputPriorityPorts_3_4; // @[Mux.scala 19:72:@11739.4]
  wire  inputPriorityPorts_3_5; // @[Mux.scala 19:72:@11741.4]
  wire  inputPriorityPorts_3_6; // @[Mux.scala 19:72:@11743.4]
  wire  inputPriorityPorts_3_7; // @[Mux.scala 19:72:@11745.4]
  wire [7:0] _T_29932; // @[Mux.scala 31:69:@11775.4]
  wire [7:0] _T_29933; // @[Mux.scala 31:69:@11776.4]
  wire [7:0] _T_29934; // @[Mux.scala 31:69:@11777.4]
  wire [7:0] _T_29935; // @[Mux.scala 31:69:@11778.4]
  wire [7:0] _T_29936; // @[Mux.scala 31:69:@11779.4]
  wire [7:0] _T_29937; // @[Mux.scala 31:69:@11780.4]
  wire [7:0] _T_29938; // @[Mux.scala 31:69:@11781.4]
  wire [7:0] _T_29939; // @[Mux.scala 31:69:@11782.4]
  wire  _T_29940; // @[OneHot.scala 66:30:@11783.4]
  wire  _T_29941; // @[OneHot.scala 66:30:@11784.4]
  wire  _T_29942; // @[OneHot.scala 66:30:@11785.4]
  wire  _T_29943; // @[OneHot.scala 66:30:@11786.4]
  wire  _T_29944; // @[OneHot.scala 66:30:@11787.4]
  wire  _T_29945; // @[OneHot.scala 66:30:@11788.4]
  wire  _T_29946; // @[OneHot.scala 66:30:@11789.4]
  wire  _T_29947; // @[OneHot.scala 66:30:@11790.4]
  wire [7:0] _T_29972; // @[Mux.scala 31:69:@11800.4]
  wire [7:0] _T_29973; // @[Mux.scala 31:69:@11801.4]
  wire [7:0] _T_29974; // @[Mux.scala 31:69:@11802.4]
  wire [7:0] _T_29975; // @[Mux.scala 31:69:@11803.4]
  wire [7:0] _T_29976; // @[Mux.scala 31:69:@11804.4]
  wire [7:0] _T_29977; // @[Mux.scala 31:69:@11805.4]
  wire [7:0] _T_29978; // @[Mux.scala 31:69:@11806.4]
  wire [7:0] _T_29979; // @[Mux.scala 31:69:@11807.4]
  wire  _T_29980; // @[OneHot.scala 66:30:@11808.4]
  wire  _T_29981; // @[OneHot.scala 66:30:@11809.4]
  wire  _T_29982; // @[OneHot.scala 66:30:@11810.4]
  wire  _T_29983; // @[OneHot.scala 66:30:@11811.4]
  wire  _T_29984; // @[OneHot.scala 66:30:@11812.4]
  wire  _T_29985; // @[OneHot.scala 66:30:@11813.4]
  wire  _T_29986; // @[OneHot.scala 66:30:@11814.4]
  wire  _T_29987; // @[OneHot.scala 66:30:@11815.4]
  wire [7:0] _T_30012; // @[Mux.scala 31:69:@11825.4]
  wire [7:0] _T_30013; // @[Mux.scala 31:69:@11826.4]
  wire [7:0] _T_30014; // @[Mux.scala 31:69:@11827.4]
  wire [7:0] _T_30015; // @[Mux.scala 31:69:@11828.4]
  wire [7:0] _T_30016; // @[Mux.scala 31:69:@11829.4]
  wire [7:0] _T_30017; // @[Mux.scala 31:69:@11830.4]
  wire [7:0] _T_30018; // @[Mux.scala 31:69:@11831.4]
  wire [7:0] _T_30019; // @[Mux.scala 31:69:@11832.4]
  wire  _T_30020; // @[OneHot.scala 66:30:@11833.4]
  wire  _T_30021; // @[OneHot.scala 66:30:@11834.4]
  wire  _T_30022; // @[OneHot.scala 66:30:@11835.4]
  wire  _T_30023; // @[OneHot.scala 66:30:@11836.4]
  wire  _T_30024; // @[OneHot.scala 66:30:@11837.4]
  wire  _T_30025; // @[OneHot.scala 66:30:@11838.4]
  wire  _T_30026; // @[OneHot.scala 66:30:@11839.4]
  wire  _T_30027; // @[OneHot.scala 66:30:@11840.4]
  wire [7:0] _T_30052; // @[Mux.scala 31:69:@11850.4]
  wire [7:0] _T_30053; // @[Mux.scala 31:69:@11851.4]
  wire [7:0] _T_30054; // @[Mux.scala 31:69:@11852.4]
  wire [7:0] _T_30055; // @[Mux.scala 31:69:@11853.4]
  wire [7:0] _T_30056; // @[Mux.scala 31:69:@11854.4]
  wire [7:0] _T_30057; // @[Mux.scala 31:69:@11855.4]
  wire [7:0] _T_30058; // @[Mux.scala 31:69:@11856.4]
  wire [7:0] _T_30059; // @[Mux.scala 31:69:@11857.4]
  wire  _T_30060; // @[OneHot.scala 66:30:@11858.4]
  wire  _T_30061; // @[OneHot.scala 66:30:@11859.4]
  wire  _T_30062; // @[OneHot.scala 66:30:@11860.4]
  wire  _T_30063; // @[OneHot.scala 66:30:@11861.4]
  wire  _T_30064; // @[OneHot.scala 66:30:@11862.4]
  wire  _T_30065; // @[OneHot.scala 66:30:@11863.4]
  wire  _T_30066; // @[OneHot.scala 66:30:@11864.4]
  wire  _T_30067; // @[OneHot.scala 66:30:@11865.4]
  wire [7:0] _T_30092; // @[Mux.scala 31:69:@11875.4]
  wire [7:0] _T_30093; // @[Mux.scala 31:69:@11876.4]
  wire [7:0] _T_30094; // @[Mux.scala 31:69:@11877.4]
  wire [7:0] _T_30095; // @[Mux.scala 31:69:@11878.4]
  wire [7:0] _T_30096; // @[Mux.scala 31:69:@11879.4]
  wire [7:0] _T_30097; // @[Mux.scala 31:69:@11880.4]
  wire [7:0] _T_30098; // @[Mux.scala 31:69:@11881.4]
  wire [7:0] _T_30099; // @[Mux.scala 31:69:@11882.4]
  wire  _T_30100; // @[OneHot.scala 66:30:@11883.4]
  wire  _T_30101; // @[OneHot.scala 66:30:@11884.4]
  wire  _T_30102; // @[OneHot.scala 66:30:@11885.4]
  wire  _T_30103; // @[OneHot.scala 66:30:@11886.4]
  wire  _T_30104; // @[OneHot.scala 66:30:@11887.4]
  wire  _T_30105; // @[OneHot.scala 66:30:@11888.4]
  wire  _T_30106; // @[OneHot.scala 66:30:@11889.4]
  wire  _T_30107; // @[OneHot.scala 66:30:@11890.4]
  wire [7:0] _T_30132; // @[Mux.scala 31:69:@11900.4]
  wire [7:0] _T_30133; // @[Mux.scala 31:69:@11901.4]
  wire [7:0] _T_30134; // @[Mux.scala 31:69:@11902.4]
  wire [7:0] _T_30135; // @[Mux.scala 31:69:@11903.4]
  wire [7:0] _T_30136; // @[Mux.scala 31:69:@11904.4]
  wire [7:0] _T_30137; // @[Mux.scala 31:69:@11905.4]
  wire [7:0] _T_30138; // @[Mux.scala 31:69:@11906.4]
  wire [7:0] _T_30139; // @[Mux.scala 31:69:@11907.4]
  wire  _T_30140; // @[OneHot.scala 66:30:@11908.4]
  wire  _T_30141; // @[OneHot.scala 66:30:@11909.4]
  wire  _T_30142; // @[OneHot.scala 66:30:@11910.4]
  wire  _T_30143; // @[OneHot.scala 66:30:@11911.4]
  wire  _T_30144; // @[OneHot.scala 66:30:@11912.4]
  wire  _T_30145; // @[OneHot.scala 66:30:@11913.4]
  wire  _T_30146; // @[OneHot.scala 66:30:@11914.4]
  wire  _T_30147; // @[OneHot.scala 66:30:@11915.4]
  wire [7:0] _T_30172; // @[Mux.scala 31:69:@11925.4]
  wire [7:0] _T_30173; // @[Mux.scala 31:69:@11926.4]
  wire [7:0] _T_30174; // @[Mux.scala 31:69:@11927.4]
  wire [7:0] _T_30175; // @[Mux.scala 31:69:@11928.4]
  wire [7:0] _T_30176; // @[Mux.scala 31:69:@11929.4]
  wire [7:0] _T_30177; // @[Mux.scala 31:69:@11930.4]
  wire [7:0] _T_30178; // @[Mux.scala 31:69:@11931.4]
  wire [7:0] _T_30179; // @[Mux.scala 31:69:@11932.4]
  wire  _T_30180; // @[OneHot.scala 66:30:@11933.4]
  wire  _T_30181; // @[OneHot.scala 66:30:@11934.4]
  wire  _T_30182; // @[OneHot.scala 66:30:@11935.4]
  wire  _T_30183; // @[OneHot.scala 66:30:@11936.4]
  wire  _T_30184; // @[OneHot.scala 66:30:@11937.4]
  wire  _T_30185; // @[OneHot.scala 66:30:@11938.4]
  wire  _T_30186; // @[OneHot.scala 66:30:@11939.4]
  wire  _T_30187; // @[OneHot.scala 66:30:@11940.4]
  wire [7:0] _T_30212; // @[Mux.scala 31:69:@11950.4]
  wire [7:0] _T_30213; // @[Mux.scala 31:69:@11951.4]
  wire [7:0] _T_30214; // @[Mux.scala 31:69:@11952.4]
  wire [7:0] _T_30215; // @[Mux.scala 31:69:@11953.4]
  wire [7:0] _T_30216; // @[Mux.scala 31:69:@11954.4]
  wire [7:0] _T_30217; // @[Mux.scala 31:69:@11955.4]
  wire [7:0] _T_30218; // @[Mux.scala 31:69:@11956.4]
  wire [7:0] _T_30219; // @[Mux.scala 31:69:@11957.4]
  wire  _T_30220; // @[OneHot.scala 66:30:@11958.4]
  wire  _T_30221; // @[OneHot.scala 66:30:@11959.4]
  wire  _T_30222; // @[OneHot.scala 66:30:@11960.4]
  wire  _T_30223; // @[OneHot.scala 66:30:@11961.4]
  wire  _T_30224; // @[OneHot.scala 66:30:@11962.4]
  wire  _T_30225; // @[OneHot.scala 66:30:@11963.4]
  wire  _T_30226; // @[OneHot.scala 66:30:@11964.4]
  wire  _T_30227; // @[OneHot.scala 66:30:@11965.4]
  wire [7:0] _T_30268; // @[Mux.scala 19:72:@11981.4]
  wire [7:0] _T_30270; // @[Mux.scala 19:72:@11982.4]
  wire [7:0] _T_30277; // @[Mux.scala 19:72:@11989.4]
  wire [7:0] _T_30279; // @[Mux.scala 19:72:@11990.4]
  wire [7:0] _T_30286; // @[Mux.scala 19:72:@11997.4]
  wire [7:0] _T_30288; // @[Mux.scala 19:72:@11998.4]
  wire [7:0] _T_30295; // @[Mux.scala 19:72:@12005.4]
  wire [7:0] _T_30297; // @[Mux.scala 19:72:@12006.4]
  wire [7:0] _T_30304; // @[Mux.scala 19:72:@12013.4]
  wire [7:0] _T_30306; // @[Mux.scala 19:72:@12014.4]
  wire [7:0] _T_30313; // @[Mux.scala 19:72:@12021.4]
  wire [7:0] _T_30315; // @[Mux.scala 19:72:@12022.4]
  wire [7:0] _T_30322; // @[Mux.scala 19:72:@12029.4]
  wire [7:0] _T_30324; // @[Mux.scala 19:72:@12030.4]
  wire [7:0] _T_30331; // @[Mux.scala 19:72:@12037.4]
  wire [7:0] _T_30333; // @[Mux.scala 19:72:@12038.4]
  wire [7:0] _T_30334; // @[Mux.scala 19:72:@12039.4]
  wire [7:0] _T_30335; // @[Mux.scala 19:72:@12040.4]
  wire [7:0] _T_30336; // @[Mux.scala 19:72:@12041.4]
  wire [7:0] _T_30337; // @[Mux.scala 19:72:@12042.4]
  wire [7:0] _T_30338; // @[Mux.scala 19:72:@12043.4]
  wire [7:0] _T_30339; // @[Mux.scala 19:72:@12044.4]
  wire [7:0] _T_30340; // @[Mux.scala 19:72:@12045.4]
  wire  outputPriorityPorts_3_0; // @[Mux.scala 19:72:@12049.4]
  wire  outputPriorityPorts_3_1; // @[Mux.scala 19:72:@12051.4]
  wire  outputPriorityPorts_3_2; // @[Mux.scala 19:72:@12053.4]
  wire  outputPriorityPorts_3_3; // @[Mux.scala 19:72:@12055.4]
  wire  outputPriorityPorts_3_4; // @[Mux.scala 19:72:@12057.4]
  wire  outputPriorityPorts_3_5; // @[Mux.scala 19:72:@12059.4]
  wire  outputPriorityPorts_3_6; // @[Mux.scala 19:72:@12061.4]
  wire  outputPriorityPorts_3_7; // @[Mux.scala 19:72:@12063.4]
  wire  _T_30420; // @[LoadQueue.scala 298:83:@12074.4]
  wire  _T_30423; // @[LoadQueue.scala 298:83:@12076.4]
  wire  _T_30426; // @[LoadQueue.scala 298:83:@12078.4]
  wire  _T_30429; // @[LoadQueue.scala 298:83:@12080.4]
  wire  _T_30432; // @[LoadQueue.scala 298:83:@12082.4]
  wire  _T_30435; // @[LoadQueue.scala 298:83:@12084.4]
  wire  _T_30438; // @[LoadQueue.scala 298:83:@12086.4]
  wire  _T_30441; // @[LoadQueue.scala 298:83:@12088.4]
  wire [7:0] _T_30492; // @[Mux.scala 31:69:@12118.4]
  wire [7:0] _T_30493; // @[Mux.scala 31:69:@12119.4]
  wire [7:0] _T_30494; // @[Mux.scala 31:69:@12120.4]
  wire [7:0] _T_30495; // @[Mux.scala 31:69:@12121.4]
  wire [7:0] _T_30496; // @[Mux.scala 31:69:@12122.4]
  wire [7:0] _T_30497; // @[Mux.scala 31:69:@12123.4]
  wire [7:0] _T_30498; // @[Mux.scala 31:69:@12124.4]
  wire [7:0] _T_30499; // @[Mux.scala 31:69:@12125.4]
  wire  _T_30500; // @[OneHot.scala 66:30:@12126.4]
  wire  _T_30501; // @[OneHot.scala 66:30:@12127.4]
  wire  _T_30502; // @[OneHot.scala 66:30:@12128.4]
  wire  _T_30503; // @[OneHot.scala 66:30:@12129.4]
  wire  _T_30504; // @[OneHot.scala 66:30:@12130.4]
  wire  _T_30505; // @[OneHot.scala 66:30:@12131.4]
  wire  _T_30506; // @[OneHot.scala 66:30:@12132.4]
  wire  _T_30507; // @[OneHot.scala 66:30:@12133.4]
  wire [7:0] _T_30532; // @[Mux.scala 31:69:@12143.4]
  wire [7:0] _T_30533; // @[Mux.scala 31:69:@12144.4]
  wire [7:0] _T_30534; // @[Mux.scala 31:69:@12145.4]
  wire [7:0] _T_30535; // @[Mux.scala 31:69:@12146.4]
  wire [7:0] _T_30536; // @[Mux.scala 31:69:@12147.4]
  wire [7:0] _T_30537; // @[Mux.scala 31:69:@12148.4]
  wire [7:0] _T_30538; // @[Mux.scala 31:69:@12149.4]
  wire [7:0] _T_30539; // @[Mux.scala 31:69:@12150.4]
  wire  _T_30540; // @[OneHot.scala 66:30:@12151.4]
  wire  _T_30541; // @[OneHot.scala 66:30:@12152.4]
  wire  _T_30542; // @[OneHot.scala 66:30:@12153.4]
  wire  _T_30543; // @[OneHot.scala 66:30:@12154.4]
  wire  _T_30544; // @[OneHot.scala 66:30:@12155.4]
  wire  _T_30545; // @[OneHot.scala 66:30:@12156.4]
  wire  _T_30546; // @[OneHot.scala 66:30:@12157.4]
  wire  _T_30547; // @[OneHot.scala 66:30:@12158.4]
  wire [7:0] _T_30572; // @[Mux.scala 31:69:@12168.4]
  wire [7:0] _T_30573; // @[Mux.scala 31:69:@12169.4]
  wire [7:0] _T_30574; // @[Mux.scala 31:69:@12170.4]
  wire [7:0] _T_30575; // @[Mux.scala 31:69:@12171.4]
  wire [7:0] _T_30576; // @[Mux.scala 31:69:@12172.4]
  wire [7:0] _T_30577; // @[Mux.scala 31:69:@12173.4]
  wire [7:0] _T_30578; // @[Mux.scala 31:69:@12174.4]
  wire [7:0] _T_30579; // @[Mux.scala 31:69:@12175.4]
  wire  _T_30580; // @[OneHot.scala 66:30:@12176.4]
  wire  _T_30581; // @[OneHot.scala 66:30:@12177.4]
  wire  _T_30582; // @[OneHot.scala 66:30:@12178.4]
  wire  _T_30583; // @[OneHot.scala 66:30:@12179.4]
  wire  _T_30584; // @[OneHot.scala 66:30:@12180.4]
  wire  _T_30585; // @[OneHot.scala 66:30:@12181.4]
  wire  _T_30586; // @[OneHot.scala 66:30:@12182.4]
  wire  _T_30587; // @[OneHot.scala 66:30:@12183.4]
  wire [7:0] _T_30612; // @[Mux.scala 31:69:@12193.4]
  wire [7:0] _T_30613; // @[Mux.scala 31:69:@12194.4]
  wire [7:0] _T_30614; // @[Mux.scala 31:69:@12195.4]
  wire [7:0] _T_30615; // @[Mux.scala 31:69:@12196.4]
  wire [7:0] _T_30616; // @[Mux.scala 31:69:@12197.4]
  wire [7:0] _T_30617; // @[Mux.scala 31:69:@12198.4]
  wire [7:0] _T_30618; // @[Mux.scala 31:69:@12199.4]
  wire [7:0] _T_30619; // @[Mux.scala 31:69:@12200.4]
  wire  _T_30620; // @[OneHot.scala 66:30:@12201.4]
  wire  _T_30621; // @[OneHot.scala 66:30:@12202.4]
  wire  _T_30622; // @[OneHot.scala 66:30:@12203.4]
  wire  _T_30623; // @[OneHot.scala 66:30:@12204.4]
  wire  _T_30624; // @[OneHot.scala 66:30:@12205.4]
  wire  _T_30625; // @[OneHot.scala 66:30:@12206.4]
  wire  _T_30626; // @[OneHot.scala 66:30:@12207.4]
  wire  _T_30627; // @[OneHot.scala 66:30:@12208.4]
  wire [7:0] _T_30652; // @[Mux.scala 31:69:@12218.4]
  wire [7:0] _T_30653; // @[Mux.scala 31:69:@12219.4]
  wire [7:0] _T_30654; // @[Mux.scala 31:69:@12220.4]
  wire [7:0] _T_30655; // @[Mux.scala 31:69:@12221.4]
  wire [7:0] _T_30656; // @[Mux.scala 31:69:@12222.4]
  wire [7:0] _T_30657; // @[Mux.scala 31:69:@12223.4]
  wire [7:0] _T_30658; // @[Mux.scala 31:69:@12224.4]
  wire [7:0] _T_30659; // @[Mux.scala 31:69:@12225.4]
  wire  _T_30660; // @[OneHot.scala 66:30:@12226.4]
  wire  _T_30661; // @[OneHot.scala 66:30:@12227.4]
  wire  _T_30662; // @[OneHot.scala 66:30:@12228.4]
  wire  _T_30663; // @[OneHot.scala 66:30:@12229.4]
  wire  _T_30664; // @[OneHot.scala 66:30:@12230.4]
  wire  _T_30665; // @[OneHot.scala 66:30:@12231.4]
  wire  _T_30666; // @[OneHot.scala 66:30:@12232.4]
  wire  _T_30667; // @[OneHot.scala 66:30:@12233.4]
  wire [7:0] _T_30692; // @[Mux.scala 31:69:@12243.4]
  wire [7:0] _T_30693; // @[Mux.scala 31:69:@12244.4]
  wire [7:0] _T_30694; // @[Mux.scala 31:69:@12245.4]
  wire [7:0] _T_30695; // @[Mux.scala 31:69:@12246.4]
  wire [7:0] _T_30696; // @[Mux.scala 31:69:@12247.4]
  wire [7:0] _T_30697; // @[Mux.scala 31:69:@12248.4]
  wire [7:0] _T_30698; // @[Mux.scala 31:69:@12249.4]
  wire [7:0] _T_30699; // @[Mux.scala 31:69:@12250.4]
  wire  _T_30700; // @[OneHot.scala 66:30:@12251.4]
  wire  _T_30701; // @[OneHot.scala 66:30:@12252.4]
  wire  _T_30702; // @[OneHot.scala 66:30:@12253.4]
  wire  _T_30703; // @[OneHot.scala 66:30:@12254.4]
  wire  _T_30704; // @[OneHot.scala 66:30:@12255.4]
  wire  _T_30705; // @[OneHot.scala 66:30:@12256.4]
  wire  _T_30706; // @[OneHot.scala 66:30:@12257.4]
  wire  _T_30707; // @[OneHot.scala 66:30:@12258.4]
  wire [7:0] _T_30732; // @[Mux.scala 31:69:@12268.4]
  wire [7:0] _T_30733; // @[Mux.scala 31:69:@12269.4]
  wire [7:0] _T_30734; // @[Mux.scala 31:69:@12270.4]
  wire [7:0] _T_30735; // @[Mux.scala 31:69:@12271.4]
  wire [7:0] _T_30736; // @[Mux.scala 31:69:@12272.4]
  wire [7:0] _T_30737; // @[Mux.scala 31:69:@12273.4]
  wire [7:0] _T_30738; // @[Mux.scala 31:69:@12274.4]
  wire [7:0] _T_30739; // @[Mux.scala 31:69:@12275.4]
  wire  _T_30740; // @[OneHot.scala 66:30:@12276.4]
  wire  _T_30741; // @[OneHot.scala 66:30:@12277.4]
  wire  _T_30742; // @[OneHot.scala 66:30:@12278.4]
  wire  _T_30743; // @[OneHot.scala 66:30:@12279.4]
  wire  _T_30744; // @[OneHot.scala 66:30:@12280.4]
  wire  _T_30745; // @[OneHot.scala 66:30:@12281.4]
  wire  _T_30746; // @[OneHot.scala 66:30:@12282.4]
  wire  _T_30747; // @[OneHot.scala 66:30:@12283.4]
  wire [7:0] _T_30772; // @[Mux.scala 31:69:@12293.4]
  wire [7:0] _T_30773; // @[Mux.scala 31:69:@12294.4]
  wire [7:0] _T_30774; // @[Mux.scala 31:69:@12295.4]
  wire [7:0] _T_30775; // @[Mux.scala 31:69:@12296.4]
  wire [7:0] _T_30776; // @[Mux.scala 31:69:@12297.4]
  wire [7:0] _T_30777; // @[Mux.scala 31:69:@12298.4]
  wire [7:0] _T_30778; // @[Mux.scala 31:69:@12299.4]
  wire [7:0] _T_30779; // @[Mux.scala 31:69:@12300.4]
  wire  _T_30780; // @[OneHot.scala 66:30:@12301.4]
  wire  _T_30781; // @[OneHot.scala 66:30:@12302.4]
  wire  _T_30782; // @[OneHot.scala 66:30:@12303.4]
  wire  _T_30783; // @[OneHot.scala 66:30:@12304.4]
  wire  _T_30784; // @[OneHot.scala 66:30:@12305.4]
  wire  _T_30785; // @[OneHot.scala 66:30:@12306.4]
  wire  _T_30786; // @[OneHot.scala 66:30:@12307.4]
  wire  _T_30787; // @[OneHot.scala 66:30:@12308.4]
  wire [7:0] _T_30828; // @[Mux.scala 19:72:@12324.4]
  wire [7:0] _T_30830; // @[Mux.scala 19:72:@12325.4]
  wire [7:0] _T_30837; // @[Mux.scala 19:72:@12332.4]
  wire [7:0] _T_30839; // @[Mux.scala 19:72:@12333.4]
  wire [7:0] _T_30846; // @[Mux.scala 19:72:@12340.4]
  wire [7:0] _T_30848; // @[Mux.scala 19:72:@12341.4]
  wire [7:0] _T_30855; // @[Mux.scala 19:72:@12348.4]
  wire [7:0] _T_30857; // @[Mux.scala 19:72:@12349.4]
  wire [7:0] _T_30864; // @[Mux.scala 19:72:@12356.4]
  wire [7:0] _T_30866; // @[Mux.scala 19:72:@12357.4]
  wire [7:0] _T_30873; // @[Mux.scala 19:72:@12364.4]
  wire [7:0] _T_30875; // @[Mux.scala 19:72:@12365.4]
  wire [7:0] _T_30882; // @[Mux.scala 19:72:@12372.4]
  wire [7:0] _T_30884; // @[Mux.scala 19:72:@12373.4]
  wire [7:0] _T_30891; // @[Mux.scala 19:72:@12380.4]
  wire [7:0] _T_30893; // @[Mux.scala 19:72:@12381.4]
  wire [7:0] _T_30894; // @[Mux.scala 19:72:@12382.4]
  wire [7:0] _T_30895; // @[Mux.scala 19:72:@12383.4]
  wire [7:0] _T_30896; // @[Mux.scala 19:72:@12384.4]
  wire [7:0] _T_30897; // @[Mux.scala 19:72:@12385.4]
  wire [7:0] _T_30898; // @[Mux.scala 19:72:@12386.4]
  wire [7:0] _T_30899; // @[Mux.scala 19:72:@12387.4]
  wire [7:0] _T_30900; // @[Mux.scala 19:72:@12388.4]
  wire  inputPriorityPorts_4_0; // @[Mux.scala 19:72:@12392.4]
  wire  inputPriorityPorts_4_1; // @[Mux.scala 19:72:@12394.4]
  wire  inputPriorityPorts_4_2; // @[Mux.scala 19:72:@12396.4]
  wire  inputPriorityPorts_4_3; // @[Mux.scala 19:72:@12398.4]
  wire  inputPriorityPorts_4_4; // @[Mux.scala 19:72:@12400.4]
  wire  inputPriorityPorts_4_5; // @[Mux.scala 19:72:@12402.4]
  wire  inputPriorityPorts_4_6; // @[Mux.scala 19:72:@12404.4]
  wire  inputPriorityPorts_4_7; // @[Mux.scala 19:72:@12406.4]
  wire [7:0] _T_31014; // @[Mux.scala 31:69:@12436.4]
  wire [7:0] _T_31015; // @[Mux.scala 31:69:@12437.4]
  wire [7:0] _T_31016; // @[Mux.scala 31:69:@12438.4]
  wire [7:0] _T_31017; // @[Mux.scala 31:69:@12439.4]
  wire [7:0] _T_31018; // @[Mux.scala 31:69:@12440.4]
  wire [7:0] _T_31019; // @[Mux.scala 31:69:@12441.4]
  wire [7:0] _T_31020; // @[Mux.scala 31:69:@12442.4]
  wire [7:0] _T_31021; // @[Mux.scala 31:69:@12443.4]
  wire  _T_31022; // @[OneHot.scala 66:30:@12444.4]
  wire  _T_31023; // @[OneHot.scala 66:30:@12445.4]
  wire  _T_31024; // @[OneHot.scala 66:30:@12446.4]
  wire  _T_31025; // @[OneHot.scala 66:30:@12447.4]
  wire  _T_31026; // @[OneHot.scala 66:30:@12448.4]
  wire  _T_31027; // @[OneHot.scala 66:30:@12449.4]
  wire  _T_31028; // @[OneHot.scala 66:30:@12450.4]
  wire  _T_31029; // @[OneHot.scala 66:30:@12451.4]
  wire [7:0] _T_31054; // @[Mux.scala 31:69:@12461.4]
  wire [7:0] _T_31055; // @[Mux.scala 31:69:@12462.4]
  wire [7:0] _T_31056; // @[Mux.scala 31:69:@12463.4]
  wire [7:0] _T_31057; // @[Mux.scala 31:69:@12464.4]
  wire [7:0] _T_31058; // @[Mux.scala 31:69:@12465.4]
  wire [7:0] _T_31059; // @[Mux.scala 31:69:@12466.4]
  wire [7:0] _T_31060; // @[Mux.scala 31:69:@12467.4]
  wire [7:0] _T_31061; // @[Mux.scala 31:69:@12468.4]
  wire  _T_31062; // @[OneHot.scala 66:30:@12469.4]
  wire  _T_31063; // @[OneHot.scala 66:30:@12470.4]
  wire  _T_31064; // @[OneHot.scala 66:30:@12471.4]
  wire  _T_31065; // @[OneHot.scala 66:30:@12472.4]
  wire  _T_31066; // @[OneHot.scala 66:30:@12473.4]
  wire  _T_31067; // @[OneHot.scala 66:30:@12474.4]
  wire  _T_31068; // @[OneHot.scala 66:30:@12475.4]
  wire  _T_31069; // @[OneHot.scala 66:30:@12476.4]
  wire [7:0] _T_31094; // @[Mux.scala 31:69:@12486.4]
  wire [7:0] _T_31095; // @[Mux.scala 31:69:@12487.4]
  wire [7:0] _T_31096; // @[Mux.scala 31:69:@12488.4]
  wire [7:0] _T_31097; // @[Mux.scala 31:69:@12489.4]
  wire [7:0] _T_31098; // @[Mux.scala 31:69:@12490.4]
  wire [7:0] _T_31099; // @[Mux.scala 31:69:@12491.4]
  wire [7:0] _T_31100; // @[Mux.scala 31:69:@12492.4]
  wire [7:0] _T_31101; // @[Mux.scala 31:69:@12493.4]
  wire  _T_31102; // @[OneHot.scala 66:30:@12494.4]
  wire  _T_31103; // @[OneHot.scala 66:30:@12495.4]
  wire  _T_31104; // @[OneHot.scala 66:30:@12496.4]
  wire  _T_31105; // @[OneHot.scala 66:30:@12497.4]
  wire  _T_31106; // @[OneHot.scala 66:30:@12498.4]
  wire  _T_31107; // @[OneHot.scala 66:30:@12499.4]
  wire  _T_31108; // @[OneHot.scala 66:30:@12500.4]
  wire  _T_31109; // @[OneHot.scala 66:30:@12501.4]
  wire [7:0] _T_31134; // @[Mux.scala 31:69:@12511.4]
  wire [7:0] _T_31135; // @[Mux.scala 31:69:@12512.4]
  wire [7:0] _T_31136; // @[Mux.scala 31:69:@12513.4]
  wire [7:0] _T_31137; // @[Mux.scala 31:69:@12514.4]
  wire [7:0] _T_31138; // @[Mux.scala 31:69:@12515.4]
  wire [7:0] _T_31139; // @[Mux.scala 31:69:@12516.4]
  wire [7:0] _T_31140; // @[Mux.scala 31:69:@12517.4]
  wire [7:0] _T_31141; // @[Mux.scala 31:69:@12518.4]
  wire  _T_31142; // @[OneHot.scala 66:30:@12519.4]
  wire  _T_31143; // @[OneHot.scala 66:30:@12520.4]
  wire  _T_31144; // @[OneHot.scala 66:30:@12521.4]
  wire  _T_31145; // @[OneHot.scala 66:30:@12522.4]
  wire  _T_31146; // @[OneHot.scala 66:30:@12523.4]
  wire  _T_31147; // @[OneHot.scala 66:30:@12524.4]
  wire  _T_31148; // @[OneHot.scala 66:30:@12525.4]
  wire  _T_31149; // @[OneHot.scala 66:30:@12526.4]
  wire [7:0] _T_31174; // @[Mux.scala 31:69:@12536.4]
  wire [7:0] _T_31175; // @[Mux.scala 31:69:@12537.4]
  wire [7:0] _T_31176; // @[Mux.scala 31:69:@12538.4]
  wire [7:0] _T_31177; // @[Mux.scala 31:69:@12539.4]
  wire [7:0] _T_31178; // @[Mux.scala 31:69:@12540.4]
  wire [7:0] _T_31179; // @[Mux.scala 31:69:@12541.4]
  wire [7:0] _T_31180; // @[Mux.scala 31:69:@12542.4]
  wire [7:0] _T_31181; // @[Mux.scala 31:69:@12543.4]
  wire  _T_31182; // @[OneHot.scala 66:30:@12544.4]
  wire  _T_31183; // @[OneHot.scala 66:30:@12545.4]
  wire  _T_31184; // @[OneHot.scala 66:30:@12546.4]
  wire  _T_31185; // @[OneHot.scala 66:30:@12547.4]
  wire  _T_31186; // @[OneHot.scala 66:30:@12548.4]
  wire  _T_31187; // @[OneHot.scala 66:30:@12549.4]
  wire  _T_31188; // @[OneHot.scala 66:30:@12550.4]
  wire  _T_31189; // @[OneHot.scala 66:30:@12551.4]
  wire [7:0] _T_31214; // @[Mux.scala 31:69:@12561.4]
  wire [7:0] _T_31215; // @[Mux.scala 31:69:@12562.4]
  wire [7:0] _T_31216; // @[Mux.scala 31:69:@12563.4]
  wire [7:0] _T_31217; // @[Mux.scala 31:69:@12564.4]
  wire [7:0] _T_31218; // @[Mux.scala 31:69:@12565.4]
  wire [7:0] _T_31219; // @[Mux.scala 31:69:@12566.4]
  wire [7:0] _T_31220; // @[Mux.scala 31:69:@12567.4]
  wire [7:0] _T_31221; // @[Mux.scala 31:69:@12568.4]
  wire  _T_31222; // @[OneHot.scala 66:30:@12569.4]
  wire  _T_31223; // @[OneHot.scala 66:30:@12570.4]
  wire  _T_31224; // @[OneHot.scala 66:30:@12571.4]
  wire  _T_31225; // @[OneHot.scala 66:30:@12572.4]
  wire  _T_31226; // @[OneHot.scala 66:30:@12573.4]
  wire  _T_31227; // @[OneHot.scala 66:30:@12574.4]
  wire  _T_31228; // @[OneHot.scala 66:30:@12575.4]
  wire  _T_31229; // @[OneHot.scala 66:30:@12576.4]
  wire [7:0] _T_31254; // @[Mux.scala 31:69:@12586.4]
  wire [7:0] _T_31255; // @[Mux.scala 31:69:@12587.4]
  wire [7:0] _T_31256; // @[Mux.scala 31:69:@12588.4]
  wire [7:0] _T_31257; // @[Mux.scala 31:69:@12589.4]
  wire [7:0] _T_31258; // @[Mux.scala 31:69:@12590.4]
  wire [7:0] _T_31259; // @[Mux.scala 31:69:@12591.4]
  wire [7:0] _T_31260; // @[Mux.scala 31:69:@12592.4]
  wire [7:0] _T_31261; // @[Mux.scala 31:69:@12593.4]
  wire  _T_31262; // @[OneHot.scala 66:30:@12594.4]
  wire  _T_31263; // @[OneHot.scala 66:30:@12595.4]
  wire  _T_31264; // @[OneHot.scala 66:30:@12596.4]
  wire  _T_31265; // @[OneHot.scala 66:30:@12597.4]
  wire  _T_31266; // @[OneHot.scala 66:30:@12598.4]
  wire  _T_31267; // @[OneHot.scala 66:30:@12599.4]
  wire  _T_31268; // @[OneHot.scala 66:30:@12600.4]
  wire  _T_31269; // @[OneHot.scala 66:30:@12601.4]
  wire [7:0] _T_31294; // @[Mux.scala 31:69:@12611.4]
  wire [7:0] _T_31295; // @[Mux.scala 31:69:@12612.4]
  wire [7:0] _T_31296; // @[Mux.scala 31:69:@12613.4]
  wire [7:0] _T_31297; // @[Mux.scala 31:69:@12614.4]
  wire [7:0] _T_31298; // @[Mux.scala 31:69:@12615.4]
  wire [7:0] _T_31299; // @[Mux.scala 31:69:@12616.4]
  wire [7:0] _T_31300; // @[Mux.scala 31:69:@12617.4]
  wire [7:0] _T_31301; // @[Mux.scala 31:69:@12618.4]
  wire  _T_31302; // @[OneHot.scala 66:30:@12619.4]
  wire  _T_31303; // @[OneHot.scala 66:30:@12620.4]
  wire  _T_31304; // @[OneHot.scala 66:30:@12621.4]
  wire  _T_31305; // @[OneHot.scala 66:30:@12622.4]
  wire  _T_31306; // @[OneHot.scala 66:30:@12623.4]
  wire  _T_31307; // @[OneHot.scala 66:30:@12624.4]
  wire  _T_31308; // @[OneHot.scala 66:30:@12625.4]
  wire  _T_31309; // @[OneHot.scala 66:30:@12626.4]
  wire [7:0] _T_31350; // @[Mux.scala 19:72:@12642.4]
  wire [7:0] _T_31352; // @[Mux.scala 19:72:@12643.4]
  wire [7:0] _T_31359; // @[Mux.scala 19:72:@12650.4]
  wire [7:0] _T_31361; // @[Mux.scala 19:72:@12651.4]
  wire [7:0] _T_31368; // @[Mux.scala 19:72:@12658.4]
  wire [7:0] _T_31370; // @[Mux.scala 19:72:@12659.4]
  wire [7:0] _T_31377; // @[Mux.scala 19:72:@12666.4]
  wire [7:0] _T_31379; // @[Mux.scala 19:72:@12667.4]
  wire [7:0] _T_31386; // @[Mux.scala 19:72:@12674.4]
  wire [7:0] _T_31388; // @[Mux.scala 19:72:@12675.4]
  wire [7:0] _T_31395; // @[Mux.scala 19:72:@12682.4]
  wire [7:0] _T_31397; // @[Mux.scala 19:72:@12683.4]
  wire [7:0] _T_31404; // @[Mux.scala 19:72:@12690.4]
  wire [7:0] _T_31406; // @[Mux.scala 19:72:@12691.4]
  wire [7:0] _T_31413; // @[Mux.scala 19:72:@12698.4]
  wire [7:0] _T_31415; // @[Mux.scala 19:72:@12699.4]
  wire [7:0] _T_31416; // @[Mux.scala 19:72:@12700.4]
  wire [7:0] _T_31417; // @[Mux.scala 19:72:@12701.4]
  wire [7:0] _T_31418; // @[Mux.scala 19:72:@12702.4]
  wire [7:0] _T_31419; // @[Mux.scala 19:72:@12703.4]
  wire [7:0] _T_31420; // @[Mux.scala 19:72:@12704.4]
  wire [7:0] _T_31421; // @[Mux.scala 19:72:@12705.4]
  wire [7:0] _T_31422; // @[Mux.scala 19:72:@12706.4]
  wire  outputPriorityPorts_4_0; // @[Mux.scala 19:72:@12710.4]
  wire  outputPriorityPorts_4_1; // @[Mux.scala 19:72:@12712.4]
  wire  outputPriorityPorts_4_2; // @[Mux.scala 19:72:@12714.4]
  wire  outputPriorityPorts_4_3; // @[Mux.scala 19:72:@12716.4]
  wire  outputPriorityPorts_4_4; // @[Mux.scala 19:72:@12718.4]
  wire  outputPriorityPorts_4_5; // @[Mux.scala 19:72:@12720.4]
  wire  outputPriorityPorts_4_6; // @[Mux.scala 19:72:@12722.4]
  wire  outputPriorityPorts_4_7; // @[Mux.scala 19:72:@12724.4]
  wire  _T_31501; // @[LoadQueue.scala 313:47:@12738.6]
  wire  _T_31502; // @[LoadQueue.scala 313:47:@12739.6]
  wire  _T_31503; // @[LoadQueue.scala 313:47:@12740.6]
  wire  _T_31504; // @[LoadQueue.scala 313:47:@12741.6]
  wire  _T_31505; // @[LoadQueue.scala 313:47:@12742.6]
  wire  _T_31519; // @[LoadQueue.scala 314:26:@12750.6]
  wire  _T_31520; // @[LoadQueue.scala 314:26:@12751.6]
  wire  _T_31521; // @[LoadQueue.scala 314:26:@12752.6]
  wire  _T_31522; // @[LoadQueue.scala 314:26:@12753.6]
  wire [4:0] _T_31526; // @[OneHot.scala 18:45:@12758.8]
  wire  _T_31527; // @[OneHot.scala 26:18:@12759.8]
  wire [3:0] _T_31528; // @[OneHot.scala 27:18:@12760.8]
  wire [3:0] _GEN_814; // @[OneHot.scala 28:28:@12762.8]
  wire [3:0] _T_31531; // @[OneHot.scala 28:28:@12762.8]
  wire [1:0] _T_31532; // @[OneHot.scala 26:18:@12763.8]
  wire [1:0] _T_31533; // @[OneHot.scala 27:18:@12764.8]
  wire  _T_31535; // @[OneHot.scala 28:14:@12765.8]
  wire [1:0] _T_31536; // @[OneHot.scala 28:28:@12766.8]
  wire  _T_31537; // @[CircuitMath.scala 30:8:@12767.8]
  wire [2:0] _T_31539; // @[Cat.scala 30:58:@12769.8]
  wire [31:0] _GEN_611; // @[LoadQueue.scala 315:29:@12770.8]
  wire [31:0] _GEN_612; // @[LoadQueue.scala 315:29:@12770.8]
  wire [31:0] _GEN_613; // @[LoadQueue.scala 315:29:@12770.8]
  wire [31:0] _GEN_614; // @[LoadQueue.scala 315:29:@12770.8]
  wire [31:0] _GEN_615; // @[LoadQueue.scala 314:36:@12754.6]
  wire  _GEN_616; // @[LoadQueue.scala 314:36:@12754.6]
  wire  _GEN_617; // @[LoadQueue.scala 308:34:@12734.4]
  wire [31:0] _GEN_618; // @[LoadQueue.scala 308:34:@12734.4]
  wire  _T_31543; // @[LoadQueue.scala 313:47:@12778.6]
  wire  _T_31544; // @[LoadQueue.scala 313:47:@12779.6]
  wire  _T_31545; // @[LoadQueue.scala 313:47:@12780.6]
  wire  _T_31546; // @[LoadQueue.scala 313:47:@12781.6]
  wire  _T_31547; // @[LoadQueue.scala 313:47:@12782.6]
  wire  _T_31561; // @[LoadQueue.scala 314:26:@12790.6]
  wire  _T_31562; // @[LoadQueue.scala 314:26:@12791.6]
  wire  _T_31563; // @[LoadQueue.scala 314:26:@12792.6]
  wire  _T_31564; // @[LoadQueue.scala 314:26:@12793.6]
  wire [4:0] _T_31568; // @[OneHot.scala 18:45:@12798.8]
  wire  _T_31569; // @[OneHot.scala 26:18:@12799.8]
  wire [3:0] _T_31570; // @[OneHot.scala 27:18:@12800.8]
  wire [3:0] _GEN_815; // @[OneHot.scala 28:28:@12802.8]
  wire [3:0] _T_31573; // @[OneHot.scala 28:28:@12802.8]
  wire [1:0] _T_31574; // @[OneHot.scala 26:18:@12803.8]
  wire [1:0] _T_31575; // @[OneHot.scala 27:18:@12804.8]
  wire  _T_31577; // @[OneHot.scala 28:14:@12805.8]
  wire [1:0] _T_31578; // @[OneHot.scala 28:28:@12806.8]
  wire  _T_31579; // @[CircuitMath.scala 30:8:@12807.8]
  wire [2:0] _T_31581; // @[Cat.scala 30:58:@12809.8]
  wire [31:0] _GEN_620; // @[LoadQueue.scala 315:29:@12810.8]
  wire [31:0] _GEN_621; // @[LoadQueue.scala 315:29:@12810.8]
  wire [31:0] _GEN_622; // @[LoadQueue.scala 315:29:@12810.8]
  wire [31:0] _GEN_623; // @[LoadQueue.scala 315:29:@12810.8]
  wire [31:0] _GEN_624; // @[LoadQueue.scala 314:36:@12794.6]
  wire  _GEN_625; // @[LoadQueue.scala 314:36:@12794.6]
  wire  _GEN_626; // @[LoadQueue.scala 308:34:@12774.4]
  wire [31:0] _GEN_627; // @[LoadQueue.scala 308:34:@12774.4]
  wire  _T_31585; // @[LoadQueue.scala 313:47:@12818.6]
  wire  _T_31586; // @[LoadQueue.scala 313:47:@12819.6]
  wire  _T_31587; // @[LoadQueue.scala 313:47:@12820.6]
  wire  _T_31588; // @[LoadQueue.scala 313:47:@12821.6]
  wire  _T_31589; // @[LoadQueue.scala 313:47:@12822.6]
  wire  _T_31603; // @[LoadQueue.scala 314:26:@12830.6]
  wire  _T_31604; // @[LoadQueue.scala 314:26:@12831.6]
  wire  _T_31605; // @[LoadQueue.scala 314:26:@12832.6]
  wire  _T_31606; // @[LoadQueue.scala 314:26:@12833.6]
  wire [4:0] _T_31610; // @[OneHot.scala 18:45:@12838.8]
  wire  _T_31611; // @[OneHot.scala 26:18:@12839.8]
  wire [3:0] _T_31612; // @[OneHot.scala 27:18:@12840.8]
  wire [3:0] _GEN_816; // @[OneHot.scala 28:28:@12842.8]
  wire [3:0] _T_31615; // @[OneHot.scala 28:28:@12842.8]
  wire [1:0] _T_31616; // @[OneHot.scala 26:18:@12843.8]
  wire [1:0] _T_31617; // @[OneHot.scala 27:18:@12844.8]
  wire  _T_31619; // @[OneHot.scala 28:14:@12845.8]
  wire [1:0] _T_31620; // @[OneHot.scala 28:28:@12846.8]
  wire  _T_31621; // @[CircuitMath.scala 30:8:@12847.8]
  wire [2:0] _T_31623; // @[Cat.scala 30:58:@12849.8]
  wire [31:0] _GEN_629; // @[LoadQueue.scala 315:29:@12850.8]
  wire [31:0] _GEN_630; // @[LoadQueue.scala 315:29:@12850.8]
  wire [31:0] _GEN_631; // @[LoadQueue.scala 315:29:@12850.8]
  wire [31:0] _GEN_632; // @[LoadQueue.scala 315:29:@12850.8]
  wire [31:0] _GEN_633; // @[LoadQueue.scala 314:36:@12834.6]
  wire  _GEN_634; // @[LoadQueue.scala 314:36:@12834.6]
  wire  _GEN_635; // @[LoadQueue.scala 308:34:@12814.4]
  wire [31:0] _GEN_636; // @[LoadQueue.scala 308:34:@12814.4]
  wire  _T_31627; // @[LoadQueue.scala 313:47:@12858.6]
  wire  _T_31628; // @[LoadQueue.scala 313:47:@12859.6]
  wire  _T_31629; // @[LoadQueue.scala 313:47:@12860.6]
  wire  _T_31630; // @[LoadQueue.scala 313:47:@12861.6]
  wire  _T_31631; // @[LoadQueue.scala 313:47:@12862.6]
  wire  _T_31645; // @[LoadQueue.scala 314:26:@12870.6]
  wire  _T_31646; // @[LoadQueue.scala 314:26:@12871.6]
  wire  _T_31647; // @[LoadQueue.scala 314:26:@12872.6]
  wire  _T_31648; // @[LoadQueue.scala 314:26:@12873.6]
  wire [4:0] _T_31652; // @[OneHot.scala 18:45:@12878.8]
  wire  _T_31653; // @[OneHot.scala 26:18:@12879.8]
  wire [3:0] _T_31654; // @[OneHot.scala 27:18:@12880.8]
  wire [3:0] _GEN_817; // @[OneHot.scala 28:28:@12882.8]
  wire [3:0] _T_31657; // @[OneHot.scala 28:28:@12882.8]
  wire [1:0] _T_31658; // @[OneHot.scala 26:18:@12883.8]
  wire [1:0] _T_31659; // @[OneHot.scala 27:18:@12884.8]
  wire  _T_31661; // @[OneHot.scala 28:14:@12885.8]
  wire [1:0] _T_31662; // @[OneHot.scala 28:28:@12886.8]
  wire  _T_31663; // @[CircuitMath.scala 30:8:@12887.8]
  wire [2:0] _T_31665; // @[Cat.scala 30:58:@12889.8]
  wire [31:0] _GEN_638; // @[LoadQueue.scala 315:29:@12890.8]
  wire [31:0] _GEN_639; // @[LoadQueue.scala 315:29:@12890.8]
  wire [31:0] _GEN_640; // @[LoadQueue.scala 315:29:@12890.8]
  wire [31:0] _GEN_641; // @[LoadQueue.scala 315:29:@12890.8]
  wire [31:0] _GEN_642; // @[LoadQueue.scala 314:36:@12874.6]
  wire  _GEN_643; // @[LoadQueue.scala 314:36:@12874.6]
  wire  _GEN_644; // @[LoadQueue.scala 308:34:@12854.4]
  wire [31:0] _GEN_645; // @[LoadQueue.scala 308:34:@12854.4]
  wire  _T_31669; // @[LoadQueue.scala 313:47:@12898.6]
  wire  _T_31670; // @[LoadQueue.scala 313:47:@12899.6]
  wire  _T_31671; // @[LoadQueue.scala 313:47:@12900.6]
  wire  _T_31672; // @[LoadQueue.scala 313:47:@12901.6]
  wire  _T_31673; // @[LoadQueue.scala 313:47:@12902.6]
  wire  _T_31687; // @[LoadQueue.scala 314:26:@12910.6]
  wire  _T_31688; // @[LoadQueue.scala 314:26:@12911.6]
  wire  _T_31689; // @[LoadQueue.scala 314:26:@12912.6]
  wire  _T_31690; // @[LoadQueue.scala 314:26:@12913.6]
  wire [4:0] _T_31694; // @[OneHot.scala 18:45:@12918.8]
  wire  _T_31695; // @[OneHot.scala 26:18:@12919.8]
  wire [3:0] _T_31696; // @[OneHot.scala 27:18:@12920.8]
  wire [3:0] _GEN_818; // @[OneHot.scala 28:28:@12922.8]
  wire [3:0] _T_31699; // @[OneHot.scala 28:28:@12922.8]
  wire [1:0] _T_31700; // @[OneHot.scala 26:18:@12923.8]
  wire [1:0] _T_31701; // @[OneHot.scala 27:18:@12924.8]
  wire  _T_31703; // @[OneHot.scala 28:14:@12925.8]
  wire [1:0] _T_31704; // @[OneHot.scala 28:28:@12926.8]
  wire  _T_31705; // @[CircuitMath.scala 30:8:@12927.8]
  wire [2:0] _T_31707; // @[Cat.scala 30:58:@12929.8]
  wire [31:0] _GEN_647; // @[LoadQueue.scala 315:29:@12930.8]
  wire [31:0] _GEN_648; // @[LoadQueue.scala 315:29:@12930.8]
  wire [31:0] _GEN_649; // @[LoadQueue.scala 315:29:@12930.8]
  wire [31:0] _GEN_650; // @[LoadQueue.scala 315:29:@12930.8]
  wire [31:0] _GEN_651; // @[LoadQueue.scala 314:36:@12914.6]
  wire  _GEN_652; // @[LoadQueue.scala 314:36:@12914.6]
  wire  _GEN_653; // @[LoadQueue.scala 308:34:@12894.4]
  wire [31:0] _GEN_654; // @[LoadQueue.scala 308:34:@12894.4]
  wire  _T_31711; // @[LoadQueue.scala 313:47:@12938.6]
  wire  _T_31712; // @[LoadQueue.scala 313:47:@12939.6]
  wire  _T_31713; // @[LoadQueue.scala 313:47:@12940.6]
  wire  _T_31714; // @[LoadQueue.scala 313:47:@12941.6]
  wire  _T_31715; // @[LoadQueue.scala 313:47:@12942.6]
  wire  _T_31729; // @[LoadQueue.scala 314:26:@12950.6]
  wire  _T_31730; // @[LoadQueue.scala 314:26:@12951.6]
  wire  _T_31731; // @[LoadQueue.scala 314:26:@12952.6]
  wire  _T_31732; // @[LoadQueue.scala 314:26:@12953.6]
  wire [4:0] _T_31736; // @[OneHot.scala 18:45:@12958.8]
  wire  _T_31737; // @[OneHot.scala 26:18:@12959.8]
  wire [3:0] _T_31738; // @[OneHot.scala 27:18:@12960.8]
  wire [3:0] _GEN_819; // @[OneHot.scala 28:28:@12962.8]
  wire [3:0] _T_31741; // @[OneHot.scala 28:28:@12962.8]
  wire [1:0] _T_31742; // @[OneHot.scala 26:18:@12963.8]
  wire [1:0] _T_31743; // @[OneHot.scala 27:18:@12964.8]
  wire  _T_31745; // @[OneHot.scala 28:14:@12965.8]
  wire [1:0] _T_31746; // @[OneHot.scala 28:28:@12966.8]
  wire  _T_31747; // @[CircuitMath.scala 30:8:@12967.8]
  wire [2:0] _T_31749; // @[Cat.scala 30:58:@12969.8]
  wire [31:0] _GEN_656; // @[LoadQueue.scala 315:29:@12970.8]
  wire [31:0] _GEN_657; // @[LoadQueue.scala 315:29:@12970.8]
  wire [31:0] _GEN_658; // @[LoadQueue.scala 315:29:@12970.8]
  wire [31:0] _GEN_659; // @[LoadQueue.scala 315:29:@12970.8]
  wire [31:0] _GEN_660; // @[LoadQueue.scala 314:36:@12954.6]
  wire  _GEN_661; // @[LoadQueue.scala 314:36:@12954.6]
  wire  _GEN_662; // @[LoadQueue.scala 308:34:@12934.4]
  wire [31:0] _GEN_663; // @[LoadQueue.scala 308:34:@12934.4]
  wire  _T_31753; // @[LoadQueue.scala 313:47:@12978.6]
  wire  _T_31754; // @[LoadQueue.scala 313:47:@12979.6]
  wire  _T_31755; // @[LoadQueue.scala 313:47:@12980.6]
  wire  _T_31756; // @[LoadQueue.scala 313:47:@12981.6]
  wire  _T_31757; // @[LoadQueue.scala 313:47:@12982.6]
  wire  _T_31771; // @[LoadQueue.scala 314:26:@12990.6]
  wire  _T_31772; // @[LoadQueue.scala 314:26:@12991.6]
  wire  _T_31773; // @[LoadQueue.scala 314:26:@12992.6]
  wire  _T_31774; // @[LoadQueue.scala 314:26:@12993.6]
  wire [4:0] _T_31778; // @[OneHot.scala 18:45:@12998.8]
  wire  _T_31779; // @[OneHot.scala 26:18:@12999.8]
  wire [3:0] _T_31780; // @[OneHot.scala 27:18:@13000.8]
  wire [3:0] _GEN_820; // @[OneHot.scala 28:28:@13002.8]
  wire [3:0] _T_31783; // @[OneHot.scala 28:28:@13002.8]
  wire [1:0] _T_31784; // @[OneHot.scala 26:18:@13003.8]
  wire [1:0] _T_31785; // @[OneHot.scala 27:18:@13004.8]
  wire  _T_31787; // @[OneHot.scala 28:14:@13005.8]
  wire [1:0] _T_31788; // @[OneHot.scala 28:28:@13006.8]
  wire  _T_31789; // @[CircuitMath.scala 30:8:@13007.8]
  wire [2:0] _T_31791; // @[Cat.scala 30:58:@13009.8]
  wire [31:0] _GEN_665; // @[LoadQueue.scala 315:29:@13010.8]
  wire [31:0] _GEN_666; // @[LoadQueue.scala 315:29:@13010.8]
  wire [31:0] _GEN_667; // @[LoadQueue.scala 315:29:@13010.8]
  wire [31:0] _GEN_668; // @[LoadQueue.scala 315:29:@13010.8]
  wire [31:0] _GEN_669; // @[LoadQueue.scala 314:36:@12994.6]
  wire  _GEN_670; // @[LoadQueue.scala 314:36:@12994.6]
  wire  _GEN_671; // @[LoadQueue.scala 308:34:@12974.4]
  wire [31:0] _GEN_672; // @[LoadQueue.scala 308:34:@12974.4]
  wire  _T_31795; // @[LoadQueue.scala 313:47:@13018.6]
  wire  _T_31796; // @[LoadQueue.scala 313:47:@13019.6]
  wire  _T_31797; // @[LoadQueue.scala 313:47:@13020.6]
  wire  _T_31798; // @[LoadQueue.scala 313:47:@13021.6]
  wire  _T_31799; // @[LoadQueue.scala 313:47:@13022.6]
  wire  _T_31813; // @[LoadQueue.scala 314:26:@13030.6]
  wire  _T_31814; // @[LoadQueue.scala 314:26:@13031.6]
  wire  _T_31815; // @[LoadQueue.scala 314:26:@13032.6]
  wire  _T_31816; // @[LoadQueue.scala 314:26:@13033.6]
  wire [4:0] _T_31820; // @[OneHot.scala 18:45:@13038.8]
  wire  _T_31821; // @[OneHot.scala 26:18:@13039.8]
  wire [3:0] _T_31822; // @[OneHot.scala 27:18:@13040.8]
  wire [3:0] _GEN_821; // @[OneHot.scala 28:28:@13042.8]
  wire [3:0] _T_31825; // @[OneHot.scala 28:28:@13042.8]
  wire [1:0] _T_31826; // @[OneHot.scala 26:18:@13043.8]
  wire [1:0] _T_31827; // @[OneHot.scala 27:18:@13044.8]
  wire  _T_31829; // @[OneHot.scala 28:14:@13045.8]
  wire [1:0] _T_31830; // @[OneHot.scala 28:28:@13046.8]
  wire  _T_31831; // @[CircuitMath.scala 30:8:@13047.8]
  wire [2:0] _T_31833; // @[Cat.scala 30:58:@13049.8]
  wire [31:0] _GEN_674; // @[LoadQueue.scala 315:29:@13050.8]
  wire [31:0] _GEN_675; // @[LoadQueue.scala 315:29:@13050.8]
  wire [31:0] _GEN_676; // @[LoadQueue.scala 315:29:@13050.8]
  wire [31:0] _GEN_677; // @[LoadQueue.scala 315:29:@13050.8]
  wire [31:0] _GEN_678; // @[LoadQueue.scala 314:36:@13034.6]
  wire  _GEN_679; // @[LoadQueue.scala 314:36:@13034.6]
  wire  _GEN_680; // @[LoadQueue.scala 308:34:@13014.4]
  wire [31:0] _GEN_681; // @[LoadQueue.scala 308:34:@13014.4]
  wire  _T_31849; // @[LoadQueue.scala 326:108:@13055.4]
  wire  _T_31851; // @[LoadQueue.scala 327:34:@13056.4]
  wire  _T_31852; // @[LoadQueue.scala 327:31:@13057.4]
  wire  _T_31853; // @[LoadQueue.scala 327:63:@13058.4]
  wire  _T_31854; // @[LoadQueue.scala 326:108:@13059.4]
  wire  _T_31857; // @[LoadQueue.scala 327:31:@13061.4]
  wire  _T_31858; // @[LoadQueue.scala 327:63:@13062.4]
  wire  _T_31859; // @[LoadQueue.scala 326:108:@13063.4]
  wire  _T_31862; // @[LoadQueue.scala 327:31:@13065.4]
  wire  _T_31863; // @[LoadQueue.scala 327:63:@13066.4]
  wire  _T_31864; // @[LoadQueue.scala 326:108:@13067.4]
  wire  _T_31867; // @[LoadQueue.scala 327:31:@13069.4]
  wire  _T_31868; // @[LoadQueue.scala 327:63:@13070.4]
  wire  _T_31869; // @[LoadQueue.scala 326:108:@13071.4]
  wire  _T_31872; // @[LoadQueue.scala 327:31:@13073.4]
  wire  _T_31873; // @[LoadQueue.scala 327:63:@13074.4]
  wire  _T_31887; // @[LoadQueue.scala 328:51:@13082.4]
  wire  _T_31888; // @[LoadQueue.scala 328:51:@13083.4]
  wire  _T_31889; // @[LoadQueue.scala 328:51:@13084.4]
  wire  loadCompleting_0; // @[LoadQueue.scala 328:51:@13085.4]
  wire  _T_31891; // @[LoadQueue.scala 326:108:@13087.4]
  wire  _T_31893; // @[LoadQueue.scala 327:34:@13088.4]
  wire  _T_31894; // @[LoadQueue.scala 327:31:@13089.4]
  wire  _T_31895; // @[LoadQueue.scala 327:63:@13090.4]
  wire  _T_31896; // @[LoadQueue.scala 326:108:@13091.4]
  wire  _T_31899; // @[LoadQueue.scala 327:31:@13093.4]
  wire  _T_31900; // @[LoadQueue.scala 327:63:@13094.4]
  wire  _T_31901; // @[LoadQueue.scala 326:108:@13095.4]
  wire  _T_31904; // @[LoadQueue.scala 327:31:@13097.4]
  wire  _T_31905; // @[LoadQueue.scala 327:63:@13098.4]
  wire  _T_31906; // @[LoadQueue.scala 326:108:@13099.4]
  wire  _T_31909; // @[LoadQueue.scala 327:31:@13101.4]
  wire  _T_31910; // @[LoadQueue.scala 327:63:@13102.4]
  wire  _T_31911; // @[LoadQueue.scala 326:108:@13103.4]
  wire  _T_31914; // @[LoadQueue.scala 327:31:@13105.4]
  wire  _T_31915; // @[LoadQueue.scala 327:63:@13106.4]
  wire  _T_31929; // @[LoadQueue.scala 328:51:@13114.4]
  wire  _T_31930; // @[LoadQueue.scala 328:51:@13115.4]
  wire  _T_31931; // @[LoadQueue.scala 328:51:@13116.4]
  wire  loadCompleting_1; // @[LoadQueue.scala 328:51:@13117.4]
  wire  _T_31933; // @[LoadQueue.scala 326:108:@13119.4]
  wire  _T_31935; // @[LoadQueue.scala 327:34:@13120.4]
  wire  _T_31936; // @[LoadQueue.scala 327:31:@13121.4]
  wire  _T_31937; // @[LoadQueue.scala 327:63:@13122.4]
  wire  _T_31938; // @[LoadQueue.scala 326:108:@13123.4]
  wire  _T_31941; // @[LoadQueue.scala 327:31:@13125.4]
  wire  _T_31942; // @[LoadQueue.scala 327:63:@13126.4]
  wire  _T_31943; // @[LoadQueue.scala 326:108:@13127.4]
  wire  _T_31946; // @[LoadQueue.scala 327:31:@13129.4]
  wire  _T_31947; // @[LoadQueue.scala 327:63:@13130.4]
  wire  _T_31948; // @[LoadQueue.scala 326:108:@13131.4]
  wire  _T_31951; // @[LoadQueue.scala 327:31:@13133.4]
  wire  _T_31952; // @[LoadQueue.scala 327:63:@13134.4]
  wire  _T_31953; // @[LoadQueue.scala 326:108:@13135.4]
  wire  _T_31956; // @[LoadQueue.scala 327:31:@13137.4]
  wire  _T_31957; // @[LoadQueue.scala 327:63:@13138.4]
  wire  _T_31971; // @[LoadQueue.scala 328:51:@13146.4]
  wire  _T_31972; // @[LoadQueue.scala 328:51:@13147.4]
  wire  _T_31973; // @[LoadQueue.scala 328:51:@13148.4]
  wire  loadCompleting_2; // @[LoadQueue.scala 328:51:@13149.4]
  wire  _T_31975; // @[LoadQueue.scala 326:108:@13151.4]
  wire  _T_31977; // @[LoadQueue.scala 327:34:@13152.4]
  wire  _T_31978; // @[LoadQueue.scala 327:31:@13153.4]
  wire  _T_31979; // @[LoadQueue.scala 327:63:@13154.4]
  wire  _T_31980; // @[LoadQueue.scala 326:108:@13155.4]
  wire  _T_31983; // @[LoadQueue.scala 327:31:@13157.4]
  wire  _T_31984; // @[LoadQueue.scala 327:63:@13158.4]
  wire  _T_31985; // @[LoadQueue.scala 326:108:@13159.4]
  wire  _T_31988; // @[LoadQueue.scala 327:31:@13161.4]
  wire  _T_31989; // @[LoadQueue.scala 327:63:@13162.4]
  wire  _T_31990; // @[LoadQueue.scala 326:108:@13163.4]
  wire  _T_31993; // @[LoadQueue.scala 327:31:@13165.4]
  wire  _T_31994; // @[LoadQueue.scala 327:63:@13166.4]
  wire  _T_31995; // @[LoadQueue.scala 326:108:@13167.4]
  wire  _T_31998; // @[LoadQueue.scala 327:31:@13169.4]
  wire  _T_31999; // @[LoadQueue.scala 327:63:@13170.4]
  wire  _T_32013; // @[LoadQueue.scala 328:51:@13178.4]
  wire  _T_32014; // @[LoadQueue.scala 328:51:@13179.4]
  wire  _T_32015; // @[LoadQueue.scala 328:51:@13180.4]
  wire  loadCompleting_3; // @[LoadQueue.scala 328:51:@13181.4]
  wire  _T_32017; // @[LoadQueue.scala 326:108:@13183.4]
  wire  _T_32019; // @[LoadQueue.scala 327:34:@13184.4]
  wire  _T_32020; // @[LoadQueue.scala 327:31:@13185.4]
  wire  _T_32021; // @[LoadQueue.scala 327:63:@13186.4]
  wire  _T_32022; // @[LoadQueue.scala 326:108:@13187.4]
  wire  _T_32025; // @[LoadQueue.scala 327:31:@13189.4]
  wire  _T_32026; // @[LoadQueue.scala 327:63:@13190.4]
  wire  _T_32027; // @[LoadQueue.scala 326:108:@13191.4]
  wire  _T_32030; // @[LoadQueue.scala 327:31:@13193.4]
  wire  _T_32031; // @[LoadQueue.scala 327:63:@13194.4]
  wire  _T_32032; // @[LoadQueue.scala 326:108:@13195.4]
  wire  _T_32035; // @[LoadQueue.scala 327:31:@13197.4]
  wire  _T_32036; // @[LoadQueue.scala 327:63:@13198.4]
  wire  _T_32037; // @[LoadQueue.scala 326:108:@13199.4]
  wire  _T_32040; // @[LoadQueue.scala 327:31:@13201.4]
  wire  _T_32041; // @[LoadQueue.scala 327:63:@13202.4]
  wire  _T_32055; // @[LoadQueue.scala 328:51:@13210.4]
  wire  _T_32056; // @[LoadQueue.scala 328:51:@13211.4]
  wire  _T_32057; // @[LoadQueue.scala 328:51:@13212.4]
  wire  loadCompleting_4; // @[LoadQueue.scala 328:51:@13213.4]
  wire  _T_32059; // @[LoadQueue.scala 326:108:@13215.4]
  wire  _T_32061; // @[LoadQueue.scala 327:34:@13216.4]
  wire  _T_32062; // @[LoadQueue.scala 327:31:@13217.4]
  wire  _T_32063; // @[LoadQueue.scala 327:63:@13218.4]
  wire  _T_32064; // @[LoadQueue.scala 326:108:@13219.4]
  wire  _T_32067; // @[LoadQueue.scala 327:31:@13221.4]
  wire  _T_32068; // @[LoadQueue.scala 327:63:@13222.4]
  wire  _T_32069; // @[LoadQueue.scala 326:108:@13223.4]
  wire  _T_32072; // @[LoadQueue.scala 327:31:@13225.4]
  wire  _T_32073; // @[LoadQueue.scala 327:63:@13226.4]
  wire  _T_32074; // @[LoadQueue.scala 326:108:@13227.4]
  wire  _T_32077; // @[LoadQueue.scala 327:31:@13229.4]
  wire  _T_32078; // @[LoadQueue.scala 327:63:@13230.4]
  wire  _T_32079; // @[LoadQueue.scala 326:108:@13231.4]
  wire  _T_32082; // @[LoadQueue.scala 327:31:@13233.4]
  wire  _T_32083; // @[LoadQueue.scala 327:63:@13234.4]
  wire  _T_32097; // @[LoadQueue.scala 328:51:@13242.4]
  wire  _T_32098; // @[LoadQueue.scala 328:51:@13243.4]
  wire  _T_32099; // @[LoadQueue.scala 328:51:@13244.4]
  wire  loadCompleting_5; // @[LoadQueue.scala 328:51:@13245.4]
  wire  _T_32101; // @[LoadQueue.scala 326:108:@13247.4]
  wire  _T_32103; // @[LoadQueue.scala 327:34:@13248.4]
  wire  _T_32104; // @[LoadQueue.scala 327:31:@13249.4]
  wire  _T_32105; // @[LoadQueue.scala 327:63:@13250.4]
  wire  _T_32106; // @[LoadQueue.scala 326:108:@13251.4]
  wire  _T_32109; // @[LoadQueue.scala 327:31:@13253.4]
  wire  _T_32110; // @[LoadQueue.scala 327:63:@13254.4]
  wire  _T_32111; // @[LoadQueue.scala 326:108:@13255.4]
  wire  _T_32114; // @[LoadQueue.scala 327:31:@13257.4]
  wire  _T_32115; // @[LoadQueue.scala 327:63:@13258.4]
  wire  _T_32116; // @[LoadQueue.scala 326:108:@13259.4]
  wire  _T_32119; // @[LoadQueue.scala 327:31:@13261.4]
  wire  _T_32120; // @[LoadQueue.scala 327:63:@13262.4]
  wire  _T_32121; // @[LoadQueue.scala 326:108:@13263.4]
  wire  _T_32124; // @[LoadQueue.scala 327:31:@13265.4]
  wire  _T_32125; // @[LoadQueue.scala 327:63:@13266.4]
  wire  _T_32139; // @[LoadQueue.scala 328:51:@13274.4]
  wire  _T_32140; // @[LoadQueue.scala 328:51:@13275.4]
  wire  _T_32141; // @[LoadQueue.scala 328:51:@13276.4]
  wire  loadCompleting_6; // @[LoadQueue.scala 328:51:@13277.4]
  wire  _T_32143; // @[LoadQueue.scala 326:108:@13279.4]
  wire  _T_32145; // @[LoadQueue.scala 327:34:@13280.4]
  wire  _T_32146; // @[LoadQueue.scala 327:31:@13281.4]
  wire  _T_32147; // @[LoadQueue.scala 327:63:@13282.4]
  wire  _T_32148; // @[LoadQueue.scala 326:108:@13283.4]
  wire  _T_32151; // @[LoadQueue.scala 327:31:@13285.4]
  wire  _T_32152; // @[LoadQueue.scala 327:63:@13286.4]
  wire  _T_32153; // @[LoadQueue.scala 326:108:@13287.4]
  wire  _T_32156; // @[LoadQueue.scala 327:31:@13289.4]
  wire  _T_32157; // @[LoadQueue.scala 327:63:@13290.4]
  wire  _T_32158; // @[LoadQueue.scala 326:108:@13291.4]
  wire  _T_32161; // @[LoadQueue.scala 327:31:@13293.4]
  wire  _T_32162; // @[LoadQueue.scala 327:63:@13294.4]
  wire  _T_32163; // @[LoadQueue.scala 326:108:@13295.4]
  wire  _T_32166; // @[LoadQueue.scala 327:31:@13297.4]
  wire  _T_32167; // @[LoadQueue.scala 327:63:@13298.4]
  wire  _T_32181; // @[LoadQueue.scala 328:51:@13306.4]
  wire  _T_32182; // @[LoadQueue.scala 328:51:@13307.4]
  wire  _T_32183; // @[LoadQueue.scala 328:51:@13308.4]
  wire  loadCompleting_7; // @[LoadQueue.scala 328:51:@13309.4]
  wire  _GEN_682; // @[LoadQueue.scala 337:46:@13315.6]
  wire  _GEN_683; // @[LoadQueue.scala 335:34:@13311.4]
  wire  _GEN_684; // @[LoadQueue.scala 337:46:@13322.6]
  wire  _GEN_685; // @[LoadQueue.scala 335:34:@13318.4]
  wire  _GEN_686; // @[LoadQueue.scala 337:46:@13329.6]
  wire  _GEN_687; // @[LoadQueue.scala 335:34:@13325.4]
  wire  _GEN_688; // @[LoadQueue.scala 337:46:@13336.6]
  wire  _GEN_689; // @[LoadQueue.scala 335:34:@13332.4]
  wire  _GEN_690; // @[LoadQueue.scala 337:46:@13343.6]
  wire  _GEN_691; // @[LoadQueue.scala 335:34:@13339.4]
  wire  _GEN_692; // @[LoadQueue.scala 337:46:@13350.6]
  wire  _GEN_693; // @[LoadQueue.scala 335:34:@13346.4]
  wire  _GEN_694; // @[LoadQueue.scala 337:46:@13357.6]
  wire  _GEN_695; // @[LoadQueue.scala 335:34:@13353.4]
  wire  _GEN_696; // @[LoadQueue.scala 337:46:@13364.6]
  wire  _GEN_697; // @[LoadQueue.scala 335:34:@13360.4]
  wire  _T_32249; // @[LoadQueue.scala 348:24:@13401.4]
  wire  _T_32250; // @[LoadQueue.scala 348:24:@13402.4]
  wire  _T_32251; // @[LoadQueue.scala 348:24:@13403.4]
  wire  _T_32252; // @[LoadQueue.scala 348:24:@13404.4]
  wire  _T_32253; // @[LoadQueue.scala 348:24:@13405.4]
  wire  _T_32254; // @[LoadQueue.scala 348:24:@13406.4]
  wire  _T_32255; // @[LoadQueue.scala 348:24:@13407.4]
  wire [2:0] _T_32264; // @[Mux.scala 31:69:@13409.6]
  wire [2:0] _T_32265; // @[Mux.scala 31:69:@13410.6]
  wire [2:0] _T_32266; // @[Mux.scala 31:69:@13411.6]
  wire [2:0] _T_32267; // @[Mux.scala 31:69:@13412.6]
  wire [2:0] _T_32268; // @[Mux.scala 31:69:@13413.6]
  wire [2:0] _T_32269; // @[Mux.scala 31:69:@13414.6]
  wire [2:0] _T_32270; // @[Mux.scala 31:69:@13415.6]
  wire [31:0] _GEN_699; // @[LoadQueue.scala 349:37:@13416.6]
  wire [31:0] _GEN_700; // @[LoadQueue.scala 349:37:@13416.6]
  wire [31:0] _GEN_701; // @[LoadQueue.scala 349:37:@13416.6]
  wire [31:0] _GEN_702; // @[LoadQueue.scala 349:37:@13416.6]
  wire [31:0] _GEN_703; // @[LoadQueue.scala 349:37:@13416.6]
  wire [31:0] _GEN_704; // @[LoadQueue.scala 349:37:@13416.6]
  wire [31:0] _GEN_705; // @[LoadQueue.scala 349:37:@13416.6]
  wire  _T_32325; // @[LoadQueue.scala 348:24:@13457.4]
  wire  _T_32326; // @[LoadQueue.scala 348:24:@13458.4]
  wire  _T_32327; // @[LoadQueue.scala 348:24:@13459.4]
  wire  _T_32328; // @[LoadQueue.scala 348:24:@13460.4]
  wire  _T_32329; // @[LoadQueue.scala 348:24:@13461.4]
  wire  _T_32330; // @[LoadQueue.scala 348:24:@13462.4]
  wire  _T_32331; // @[LoadQueue.scala 348:24:@13463.4]
  wire [2:0] _T_32340; // @[Mux.scala 31:69:@13465.6]
  wire [2:0] _T_32341; // @[Mux.scala 31:69:@13466.6]
  wire [2:0] _T_32342; // @[Mux.scala 31:69:@13467.6]
  wire [2:0] _T_32343; // @[Mux.scala 31:69:@13468.6]
  wire [2:0] _T_32344; // @[Mux.scala 31:69:@13469.6]
  wire [2:0] _T_32345; // @[Mux.scala 31:69:@13470.6]
  wire [2:0] _T_32346; // @[Mux.scala 31:69:@13471.6]
  wire [31:0] _GEN_709; // @[LoadQueue.scala 349:37:@13472.6]
  wire [31:0] _GEN_710; // @[LoadQueue.scala 349:37:@13472.6]
  wire [31:0] _GEN_711; // @[LoadQueue.scala 349:37:@13472.6]
  wire [31:0] _GEN_712; // @[LoadQueue.scala 349:37:@13472.6]
  wire [31:0] _GEN_713; // @[LoadQueue.scala 349:37:@13472.6]
  wire [31:0] _GEN_714; // @[LoadQueue.scala 349:37:@13472.6]
  wire [31:0] _GEN_715; // @[LoadQueue.scala 349:37:@13472.6]
  wire  _T_32401; // @[LoadQueue.scala 348:24:@13513.4]
  wire  _T_32402; // @[LoadQueue.scala 348:24:@13514.4]
  wire  _T_32403; // @[LoadQueue.scala 348:24:@13515.4]
  wire  _T_32404; // @[LoadQueue.scala 348:24:@13516.4]
  wire  _T_32405; // @[LoadQueue.scala 348:24:@13517.4]
  wire  _T_32406; // @[LoadQueue.scala 348:24:@13518.4]
  wire  _T_32407; // @[LoadQueue.scala 348:24:@13519.4]
  wire [2:0] _T_32416; // @[Mux.scala 31:69:@13521.6]
  wire [2:0] _T_32417; // @[Mux.scala 31:69:@13522.6]
  wire [2:0] _T_32418; // @[Mux.scala 31:69:@13523.6]
  wire [2:0] _T_32419; // @[Mux.scala 31:69:@13524.6]
  wire [2:0] _T_32420; // @[Mux.scala 31:69:@13525.6]
  wire [2:0] _T_32421; // @[Mux.scala 31:69:@13526.6]
  wire [2:0] _T_32422; // @[Mux.scala 31:69:@13527.6]
  wire [31:0] _GEN_719; // @[LoadQueue.scala 349:37:@13528.6]
  wire [31:0] _GEN_720; // @[LoadQueue.scala 349:37:@13528.6]
  wire [31:0] _GEN_721; // @[LoadQueue.scala 349:37:@13528.6]
  wire [31:0] _GEN_722; // @[LoadQueue.scala 349:37:@13528.6]
  wire [31:0] _GEN_723; // @[LoadQueue.scala 349:37:@13528.6]
  wire [31:0] _GEN_724; // @[LoadQueue.scala 349:37:@13528.6]
  wire [31:0] _GEN_725; // @[LoadQueue.scala 349:37:@13528.6]
  wire  _T_32477; // @[LoadQueue.scala 348:24:@13569.4]
  wire  _T_32478; // @[LoadQueue.scala 348:24:@13570.4]
  wire  _T_32479; // @[LoadQueue.scala 348:24:@13571.4]
  wire  _T_32480; // @[LoadQueue.scala 348:24:@13572.4]
  wire  _T_32481; // @[LoadQueue.scala 348:24:@13573.4]
  wire  _T_32482; // @[LoadQueue.scala 348:24:@13574.4]
  wire  _T_32483; // @[LoadQueue.scala 348:24:@13575.4]
  wire [2:0] _T_32492; // @[Mux.scala 31:69:@13577.6]
  wire [2:0] _T_32493; // @[Mux.scala 31:69:@13578.6]
  wire [2:0] _T_32494; // @[Mux.scala 31:69:@13579.6]
  wire [2:0] _T_32495; // @[Mux.scala 31:69:@13580.6]
  wire [2:0] _T_32496; // @[Mux.scala 31:69:@13581.6]
  wire [2:0] _T_32497; // @[Mux.scala 31:69:@13582.6]
  wire [2:0] _T_32498; // @[Mux.scala 31:69:@13583.6]
  wire [31:0] _GEN_729; // @[LoadQueue.scala 349:37:@13584.6]
  wire [31:0] _GEN_730; // @[LoadQueue.scala 349:37:@13584.6]
  wire [31:0] _GEN_731; // @[LoadQueue.scala 349:37:@13584.6]
  wire [31:0] _GEN_732; // @[LoadQueue.scala 349:37:@13584.6]
  wire [31:0] _GEN_733; // @[LoadQueue.scala 349:37:@13584.6]
  wire [31:0] _GEN_734; // @[LoadQueue.scala 349:37:@13584.6]
  wire [31:0] _GEN_735; // @[LoadQueue.scala 349:37:@13584.6]
  wire  _T_32553; // @[LoadQueue.scala 348:24:@13625.4]
  wire  _T_32554; // @[LoadQueue.scala 348:24:@13626.4]
  wire  _T_32555; // @[LoadQueue.scala 348:24:@13627.4]
  wire  _T_32556; // @[LoadQueue.scala 348:24:@13628.4]
  wire  _T_32557; // @[LoadQueue.scala 348:24:@13629.4]
  wire  _T_32558; // @[LoadQueue.scala 348:24:@13630.4]
  wire  _T_32559; // @[LoadQueue.scala 348:24:@13631.4]
  wire [2:0] _T_32568; // @[Mux.scala 31:69:@13633.6]
  wire [2:0] _T_32569; // @[Mux.scala 31:69:@13634.6]
  wire [2:0] _T_32570; // @[Mux.scala 31:69:@13635.6]
  wire [2:0] _T_32571; // @[Mux.scala 31:69:@13636.6]
  wire [2:0] _T_32572; // @[Mux.scala 31:69:@13637.6]
  wire [2:0] _T_32573; // @[Mux.scala 31:69:@13638.6]
  wire [2:0] _T_32574; // @[Mux.scala 31:69:@13639.6]
  wire [31:0] _GEN_739; // @[LoadQueue.scala 349:37:@13640.6]
  wire [31:0] _GEN_740; // @[LoadQueue.scala 349:37:@13640.6]
  wire [31:0] _GEN_741; // @[LoadQueue.scala 349:37:@13640.6]
  wire [31:0] _GEN_742; // @[LoadQueue.scala 349:37:@13640.6]
  wire [31:0] _GEN_743; // @[LoadQueue.scala 349:37:@13640.6]
  wire [31:0] _GEN_744; // @[LoadQueue.scala 349:37:@13640.6]
  wire [31:0] _GEN_745; // @[LoadQueue.scala 349:37:@13640.6]
  wire  _GEN_749; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_750; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_751; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_752; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_753; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_754; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_755; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_757; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_758; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_759; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_760; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_761; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_762; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _GEN_763; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _T_32585; // @[LoadQueue.scala 363:29:@13647.4]
  wire  _T_32586; // @[LoadQueue.scala 363:63:@13648.4]
  wire  _T_32588; // @[LoadQueue.scala 363:75:@13649.4]
  wire  _T_32589; // @[LoadQueue.scala 363:72:@13650.4]
  wire  _T_32590; // @[LoadQueue.scala 363:54:@13651.4]
  wire [3:0] _T_32593; // @[util.scala 10:8:@13653.6]
  wire [3:0] _GEN_144; // @[util.scala 10:14:@13654.6]
  wire [3:0] _T_32594; // @[util.scala 10:14:@13654.6]
  wire [3:0] _GEN_764; // @[LoadQueue.scala 363:91:@13652.4]
  wire [3:0] _T_32596; // @[util.scala 10:8:@13658.6]
  wire [3:0] _GEN_145; // @[util.scala 10:14:@13659.6]
  wire [3:0] _T_32597; // @[util.scala 10:14:@13659.6]
  wire [3:0] _GEN_765; // @[LoadQueue.scala 367:20:@13657.4]
  wire  _T_32599; // @[LoadQueue.scala 371:82:@13662.4]
  wire  _T_32600; // @[LoadQueue.scala 371:79:@13663.4]
  wire  _T_32602; // @[LoadQueue.scala 371:82:@13664.4]
  wire  _T_32603; // @[LoadQueue.scala 371:79:@13665.4]
  wire  _T_32605; // @[LoadQueue.scala 371:82:@13666.4]
  wire  _T_32606; // @[LoadQueue.scala 371:79:@13667.4]
  wire  _T_32608; // @[LoadQueue.scala 371:82:@13668.4]
  wire  _T_32609; // @[LoadQueue.scala 371:79:@13669.4]
  wire  _T_32611; // @[LoadQueue.scala 371:82:@13670.4]
  wire  _T_32612; // @[LoadQueue.scala 371:79:@13671.4]
  wire  _T_32614; // @[LoadQueue.scala 371:82:@13672.4]
  wire  _T_32615; // @[LoadQueue.scala 371:79:@13673.4]
  wire  _T_32617; // @[LoadQueue.scala 371:82:@13674.4]
  wire  _T_32618; // @[LoadQueue.scala 371:79:@13675.4]
  wire  _T_32620; // @[LoadQueue.scala 371:82:@13676.4]
  wire  _T_32621; // @[LoadQueue.scala 371:79:@13677.4]
  wire  _T_32638; // @[LoadQueue.scala 371:96:@13688.4]
  wire  _T_32639; // @[LoadQueue.scala 371:96:@13689.4]
  wire  _T_32640; // @[LoadQueue.scala 371:96:@13690.4]
  wire  _T_32641; // @[LoadQueue.scala 371:96:@13691.4]
  wire  _T_32642; // @[LoadQueue.scala 371:96:@13692.4]
  wire  _T_32643; // @[LoadQueue.scala 371:96:@13693.4]
  assign _GEN_766 = {{2'd0}, tail}; // @[util.scala 14:20:@2056.4]
  assign _T_1044 = 5'h8 - _GEN_766; // @[util.scala 14:20:@2056.4]
  assign _T_1045 = $unsigned(_T_1044); // @[util.scala 14:20:@2057.4]
  assign _T_1046 = _T_1045[4:0]; // @[util.scala 14:20:@2058.4]
  assign _GEN_0 = _T_1046 % 5'h8; // @[util.scala 14:25:@2059.4]
  assign _T_1047 = _GEN_0[3:0]; // @[util.scala 14:25:@2059.4]
  assign _GEN_767 = {{1'd0}, io_bbNumLoads}; // @[LoadQueue.scala 71:46:@2060.4]
  assign _T_1048 = _T_1047 < _GEN_767; // @[LoadQueue.scala 71:46:@2060.4]
  assign initBits_0 = _T_1048 & io_bbStart; // @[LoadQueue.scala 71:63:@2061.4]
  assign _T_1053 = 5'h9 - _GEN_766; // @[util.scala 14:20:@2063.4]
  assign _T_1054 = $unsigned(_T_1053); // @[util.scala 14:20:@2064.4]
  assign _T_1055 = _T_1054[4:0]; // @[util.scala 14:20:@2065.4]
  assign _GEN_8 = _T_1055 % 5'h8; // @[util.scala 14:25:@2066.4]
  assign _T_1056 = _GEN_8[3:0]; // @[util.scala 14:25:@2066.4]
  assign _T_1057 = _T_1056 < _GEN_767; // @[LoadQueue.scala 71:46:@2067.4]
  assign initBits_1 = _T_1057 & io_bbStart; // @[LoadQueue.scala 71:63:@2068.4]
  assign _T_1062 = 5'ha - _GEN_766; // @[util.scala 14:20:@2070.4]
  assign _T_1063 = $unsigned(_T_1062); // @[util.scala 14:20:@2071.4]
  assign _T_1064 = _T_1063[4:0]; // @[util.scala 14:20:@2072.4]
  assign _GEN_18 = _T_1064 % 5'h8; // @[util.scala 14:25:@2073.4]
  assign _T_1065 = _GEN_18[3:0]; // @[util.scala 14:25:@2073.4]
  assign _T_1066 = _T_1065 < _GEN_767; // @[LoadQueue.scala 71:46:@2074.4]
  assign initBits_2 = _T_1066 & io_bbStart; // @[LoadQueue.scala 71:63:@2075.4]
  assign _T_1071 = 5'hb - _GEN_766; // @[util.scala 14:20:@2077.4]
  assign _T_1072 = $unsigned(_T_1071); // @[util.scala 14:20:@2078.4]
  assign _T_1073 = _T_1072[4:0]; // @[util.scala 14:20:@2079.4]
  assign _GEN_26 = _T_1073 % 5'h8; // @[util.scala 14:25:@2080.4]
  assign _T_1074 = _GEN_26[3:0]; // @[util.scala 14:25:@2080.4]
  assign _T_1075 = _T_1074 < _GEN_767; // @[LoadQueue.scala 71:46:@2081.4]
  assign initBits_3 = _T_1075 & io_bbStart; // @[LoadQueue.scala 71:63:@2082.4]
  assign _T_1080 = 5'hc - _GEN_766; // @[util.scala 14:20:@2084.4]
  assign _T_1081 = $unsigned(_T_1080); // @[util.scala 14:20:@2085.4]
  assign _T_1082 = _T_1081[4:0]; // @[util.scala 14:20:@2086.4]
  assign _GEN_36 = _T_1082 % 5'h8; // @[util.scala 14:25:@2087.4]
  assign _T_1083 = _GEN_36[3:0]; // @[util.scala 14:25:@2087.4]
  assign _T_1084 = _T_1083 < _GEN_767; // @[LoadQueue.scala 71:46:@2088.4]
  assign initBits_4 = _T_1084 & io_bbStart; // @[LoadQueue.scala 71:63:@2089.4]
  assign _T_1089 = 5'hd - _GEN_766; // @[util.scala 14:20:@2091.4]
  assign _T_1090 = $unsigned(_T_1089); // @[util.scala 14:20:@2092.4]
  assign _T_1091 = _T_1090[4:0]; // @[util.scala 14:20:@2093.4]
  assign _GEN_44 = _T_1091 % 5'h8; // @[util.scala 14:25:@2094.4]
  assign _T_1092 = _GEN_44[3:0]; // @[util.scala 14:25:@2094.4]
  assign _T_1093 = _T_1092 < _GEN_767; // @[LoadQueue.scala 71:46:@2095.4]
  assign initBits_5 = _T_1093 & io_bbStart; // @[LoadQueue.scala 71:63:@2096.4]
  assign _T_1098 = 5'he - _GEN_766; // @[util.scala 14:20:@2098.4]
  assign _T_1099 = $unsigned(_T_1098); // @[util.scala 14:20:@2099.4]
  assign _T_1100 = _T_1099[4:0]; // @[util.scala 14:20:@2100.4]
  assign _GEN_54 = _T_1100 % 5'h8; // @[util.scala 14:25:@2101.4]
  assign _T_1101 = _GEN_54[3:0]; // @[util.scala 14:25:@2101.4]
  assign _T_1102 = _T_1101 < _GEN_767; // @[LoadQueue.scala 71:46:@2102.4]
  assign initBits_6 = _T_1102 & io_bbStart; // @[LoadQueue.scala 71:63:@2103.4]
  assign _T_1107 = 5'hf - _GEN_766; // @[util.scala 14:20:@2105.4]
  assign _T_1108 = $unsigned(_T_1107); // @[util.scala 14:20:@2106.4]
  assign _T_1109 = _T_1108[4:0]; // @[util.scala 14:20:@2107.4]
  assign _GEN_62 = _T_1109 % 5'h8; // @[util.scala 14:25:@2108.4]
  assign _T_1110 = _GEN_62[3:0]; // @[util.scala 14:25:@2108.4]
  assign _T_1111 = _T_1110 < _GEN_767; // @[LoadQueue.scala 71:46:@2109.4]
  assign initBits_7 = _T_1111 & io_bbStart; // @[LoadQueue.scala 71:63:@2110.4]
  assign _T_1126 = allocatedEntries_0 | initBits_0; // @[LoadQueue.scala 73:78:@2120.4]
  assign _T_1127 = allocatedEntries_1 | initBits_1; // @[LoadQueue.scala 73:78:@2121.4]
  assign _T_1128 = allocatedEntries_2 | initBits_2; // @[LoadQueue.scala 73:78:@2122.4]
  assign _T_1129 = allocatedEntries_3 | initBits_3; // @[LoadQueue.scala 73:78:@2123.4]
  assign _T_1130 = allocatedEntries_4 | initBits_4; // @[LoadQueue.scala 73:78:@2124.4]
  assign _T_1131 = allocatedEntries_5 | initBits_5; // @[LoadQueue.scala 73:78:@2125.4]
  assign _T_1132 = allocatedEntries_6 | initBits_6; // @[LoadQueue.scala 73:78:@2126.4]
  assign _T_1133 = allocatedEntries_7 | initBits_7; // @[LoadQueue.scala 73:78:@2127.4]
  assign _T_1156 = _T_1047[2:0]; // @[:@2151.6]
  assign _GEN_1 = 3'h1 == _T_1156 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2152.6]
  assign _GEN_2 = 3'h2 == _T_1156 ? io_bbLoadOffsets_2 : _GEN_1; // @[LoadQueue.scala 77:20:@2152.6]
  assign _GEN_3 = 3'h3 == _T_1156 ? io_bbLoadOffsets_3 : _GEN_2; // @[LoadQueue.scala 77:20:@2152.6]
  assign _GEN_4 = 3'h4 == _T_1156 ? io_bbLoadOffsets_4 : _GEN_3; // @[LoadQueue.scala 77:20:@2152.6]
  assign _GEN_5 = 3'h5 == _T_1156 ? io_bbLoadOffsets_5 : _GEN_4; // @[LoadQueue.scala 77:20:@2152.6]
  assign _GEN_6 = 3'h6 == _T_1156 ? io_bbLoadOffsets_6 : _GEN_5; // @[LoadQueue.scala 77:20:@2152.6]
  assign _GEN_7 = 3'h7 == _T_1156 ? io_bbLoadOffsets_7 : _GEN_6; // @[LoadQueue.scala 77:20:@2152.6]
  assign _GEN_9 = 3'h1 == _T_1156 ? io_bbLoadPorts_1 : io_bbLoadPorts_0; // @[LoadQueue.scala 78:18:@2159.6]
  assign _GEN_10 = 3'h2 == _T_1156 ? io_bbLoadPorts_2 : _GEN_9; // @[LoadQueue.scala 78:18:@2159.6]
  assign _GEN_11 = 3'h3 == _T_1156 ? 3'h0 : _GEN_10; // @[LoadQueue.scala 78:18:@2159.6]
  assign _GEN_12 = 3'h4 == _T_1156 ? 3'h0 : _GEN_11; // @[LoadQueue.scala 78:18:@2159.6]
  assign _GEN_13 = 3'h5 == _T_1156 ? 3'h0 : _GEN_12; // @[LoadQueue.scala 78:18:@2159.6]
  assign _GEN_14 = 3'h6 == _T_1156 ? 3'h0 : _GEN_13; // @[LoadQueue.scala 78:18:@2159.6]
  assign _GEN_15 = 3'h7 == _T_1156 ? 3'h0 : _GEN_14; // @[LoadQueue.scala 78:18:@2159.6]
  assign _GEN_16 = initBits_0 ? _GEN_7 : offsetQ_0; // @[LoadQueue.scala 76:25:@2145.4]
  assign _GEN_17 = initBits_0 ? _GEN_15 : portQ_0; // @[LoadQueue.scala 76:25:@2145.4]
  assign _T_1174 = _T_1056[2:0]; // @[:@2167.6]
  assign _GEN_19 = 3'h1 == _T_1174 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2168.6]
  assign _GEN_20 = 3'h2 == _T_1174 ? io_bbLoadOffsets_2 : _GEN_19; // @[LoadQueue.scala 77:20:@2168.6]
  assign _GEN_21 = 3'h3 == _T_1174 ? io_bbLoadOffsets_3 : _GEN_20; // @[LoadQueue.scala 77:20:@2168.6]
  assign _GEN_22 = 3'h4 == _T_1174 ? io_bbLoadOffsets_4 : _GEN_21; // @[LoadQueue.scala 77:20:@2168.6]
  assign _GEN_23 = 3'h5 == _T_1174 ? io_bbLoadOffsets_5 : _GEN_22; // @[LoadQueue.scala 77:20:@2168.6]
  assign _GEN_24 = 3'h6 == _T_1174 ? io_bbLoadOffsets_6 : _GEN_23; // @[LoadQueue.scala 77:20:@2168.6]
  assign _GEN_25 = 3'h7 == _T_1174 ? io_bbLoadOffsets_7 : _GEN_24; // @[LoadQueue.scala 77:20:@2168.6]
  assign _GEN_27 = 3'h1 == _T_1174 ? io_bbLoadPorts_1 : io_bbLoadPorts_0; // @[LoadQueue.scala 78:18:@2175.6]
  assign _GEN_28 = 3'h2 == _T_1174 ? io_bbLoadPorts_2 : _GEN_27; // @[LoadQueue.scala 78:18:@2175.6]
  assign _GEN_29 = 3'h3 == _T_1174 ? 3'h0 : _GEN_28; // @[LoadQueue.scala 78:18:@2175.6]
  assign _GEN_30 = 3'h4 == _T_1174 ? 3'h0 : _GEN_29; // @[LoadQueue.scala 78:18:@2175.6]
  assign _GEN_31 = 3'h5 == _T_1174 ? 3'h0 : _GEN_30; // @[LoadQueue.scala 78:18:@2175.6]
  assign _GEN_32 = 3'h6 == _T_1174 ? 3'h0 : _GEN_31; // @[LoadQueue.scala 78:18:@2175.6]
  assign _GEN_33 = 3'h7 == _T_1174 ? 3'h0 : _GEN_32; // @[LoadQueue.scala 78:18:@2175.6]
  assign _GEN_34 = initBits_1 ? _GEN_25 : offsetQ_1; // @[LoadQueue.scala 76:25:@2161.4]
  assign _GEN_35 = initBits_1 ? _GEN_33 : portQ_1; // @[LoadQueue.scala 76:25:@2161.4]
  assign _T_1192 = _T_1065[2:0]; // @[:@2183.6]
  assign _GEN_37 = 3'h1 == _T_1192 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2184.6]
  assign _GEN_38 = 3'h2 == _T_1192 ? io_bbLoadOffsets_2 : _GEN_37; // @[LoadQueue.scala 77:20:@2184.6]
  assign _GEN_39 = 3'h3 == _T_1192 ? io_bbLoadOffsets_3 : _GEN_38; // @[LoadQueue.scala 77:20:@2184.6]
  assign _GEN_40 = 3'h4 == _T_1192 ? io_bbLoadOffsets_4 : _GEN_39; // @[LoadQueue.scala 77:20:@2184.6]
  assign _GEN_41 = 3'h5 == _T_1192 ? io_bbLoadOffsets_5 : _GEN_40; // @[LoadQueue.scala 77:20:@2184.6]
  assign _GEN_42 = 3'h6 == _T_1192 ? io_bbLoadOffsets_6 : _GEN_41; // @[LoadQueue.scala 77:20:@2184.6]
  assign _GEN_43 = 3'h7 == _T_1192 ? io_bbLoadOffsets_7 : _GEN_42; // @[LoadQueue.scala 77:20:@2184.6]
  assign _GEN_45 = 3'h1 == _T_1192 ? io_bbLoadPorts_1 : io_bbLoadPorts_0; // @[LoadQueue.scala 78:18:@2191.6]
  assign _GEN_46 = 3'h2 == _T_1192 ? io_bbLoadPorts_2 : _GEN_45; // @[LoadQueue.scala 78:18:@2191.6]
  assign _GEN_47 = 3'h3 == _T_1192 ? 3'h0 : _GEN_46; // @[LoadQueue.scala 78:18:@2191.6]
  assign _GEN_48 = 3'h4 == _T_1192 ? 3'h0 : _GEN_47; // @[LoadQueue.scala 78:18:@2191.6]
  assign _GEN_49 = 3'h5 == _T_1192 ? 3'h0 : _GEN_48; // @[LoadQueue.scala 78:18:@2191.6]
  assign _GEN_50 = 3'h6 == _T_1192 ? 3'h0 : _GEN_49; // @[LoadQueue.scala 78:18:@2191.6]
  assign _GEN_51 = 3'h7 == _T_1192 ? 3'h0 : _GEN_50; // @[LoadQueue.scala 78:18:@2191.6]
  assign _GEN_52 = initBits_2 ? _GEN_43 : offsetQ_2; // @[LoadQueue.scala 76:25:@2177.4]
  assign _GEN_53 = initBits_2 ? _GEN_51 : portQ_2; // @[LoadQueue.scala 76:25:@2177.4]
  assign _T_1210 = _T_1074[2:0]; // @[:@2199.6]
  assign _GEN_55 = 3'h1 == _T_1210 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2200.6]
  assign _GEN_56 = 3'h2 == _T_1210 ? io_bbLoadOffsets_2 : _GEN_55; // @[LoadQueue.scala 77:20:@2200.6]
  assign _GEN_57 = 3'h3 == _T_1210 ? io_bbLoadOffsets_3 : _GEN_56; // @[LoadQueue.scala 77:20:@2200.6]
  assign _GEN_58 = 3'h4 == _T_1210 ? io_bbLoadOffsets_4 : _GEN_57; // @[LoadQueue.scala 77:20:@2200.6]
  assign _GEN_59 = 3'h5 == _T_1210 ? io_bbLoadOffsets_5 : _GEN_58; // @[LoadQueue.scala 77:20:@2200.6]
  assign _GEN_60 = 3'h6 == _T_1210 ? io_bbLoadOffsets_6 : _GEN_59; // @[LoadQueue.scala 77:20:@2200.6]
  assign _GEN_61 = 3'h7 == _T_1210 ? io_bbLoadOffsets_7 : _GEN_60; // @[LoadQueue.scala 77:20:@2200.6]
  assign _GEN_63 = 3'h1 == _T_1210 ? io_bbLoadPorts_1 : io_bbLoadPorts_0; // @[LoadQueue.scala 78:18:@2207.6]
  assign _GEN_64 = 3'h2 == _T_1210 ? io_bbLoadPorts_2 : _GEN_63; // @[LoadQueue.scala 78:18:@2207.6]
  assign _GEN_65 = 3'h3 == _T_1210 ? 3'h0 : _GEN_64; // @[LoadQueue.scala 78:18:@2207.6]
  assign _GEN_66 = 3'h4 == _T_1210 ? 3'h0 : _GEN_65; // @[LoadQueue.scala 78:18:@2207.6]
  assign _GEN_67 = 3'h5 == _T_1210 ? 3'h0 : _GEN_66; // @[LoadQueue.scala 78:18:@2207.6]
  assign _GEN_68 = 3'h6 == _T_1210 ? 3'h0 : _GEN_67; // @[LoadQueue.scala 78:18:@2207.6]
  assign _GEN_69 = 3'h7 == _T_1210 ? 3'h0 : _GEN_68; // @[LoadQueue.scala 78:18:@2207.6]
  assign _GEN_70 = initBits_3 ? _GEN_61 : offsetQ_3; // @[LoadQueue.scala 76:25:@2193.4]
  assign _GEN_71 = initBits_3 ? _GEN_69 : portQ_3; // @[LoadQueue.scala 76:25:@2193.4]
  assign _T_1228 = _T_1083[2:0]; // @[:@2215.6]
  assign _GEN_73 = 3'h1 == _T_1228 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2216.6]
  assign _GEN_74 = 3'h2 == _T_1228 ? io_bbLoadOffsets_2 : _GEN_73; // @[LoadQueue.scala 77:20:@2216.6]
  assign _GEN_75 = 3'h3 == _T_1228 ? io_bbLoadOffsets_3 : _GEN_74; // @[LoadQueue.scala 77:20:@2216.6]
  assign _GEN_76 = 3'h4 == _T_1228 ? io_bbLoadOffsets_4 : _GEN_75; // @[LoadQueue.scala 77:20:@2216.6]
  assign _GEN_77 = 3'h5 == _T_1228 ? io_bbLoadOffsets_5 : _GEN_76; // @[LoadQueue.scala 77:20:@2216.6]
  assign _GEN_78 = 3'h6 == _T_1228 ? io_bbLoadOffsets_6 : _GEN_77; // @[LoadQueue.scala 77:20:@2216.6]
  assign _GEN_79 = 3'h7 == _T_1228 ? io_bbLoadOffsets_7 : _GEN_78; // @[LoadQueue.scala 77:20:@2216.6]
  assign _GEN_81 = 3'h1 == _T_1228 ? io_bbLoadPorts_1 : io_bbLoadPorts_0; // @[LoadQueue.scala 78:18:@2223.6]
  assign _GEN_82 = 3'h2 == _T_1228 ? io_bbLoadPorts_2 : _GEN_81; // @[LoadQueue.scala 78:18:@2223.6]
  assign _GEN_83 = 3'h3 == _T_1228 ? 3'h0 : _GEN_82; // @[LoadQueue.scala 78:18:@2223.6]
  assign _GEN_84 = 3'h4 == _T_1228 ? 3'h0 : _GEN_83; // @[LoadQueue.scala 78:18:@2223.6]
  assign _GEN_85 = 3'h5 == _T_1228 ? 3'h0 : _GEN_84; // @[LoadQueue.scala 78:18:@2223.6]
  assign _GEN_86 = 3'h6 == _T_1228 ? 3'h0 : _GEN_85; // @[LoadQueue.scala 78:18:@2223.6]
  assign _GEN_87 = 3'h7 == _T_1228 ? 3'h0 : _GEN_86; // @[LoadQueue.scala 78:18:@2223.6]
  assign _GEN_88 = initBits_4 ? _GEN_79 : offsetQ_4; // @[LoadQueue.scala 76:25:@2209.4]
  assign _GEN_89 = initBits_4 ? _GEN_87 : portQ_4; // @[LoadQueue.scala 76:25:@2209.4]
  assign _T_1246 = _T_1092[2:0]; // @[:@2231.6]
  assign _GEN_91 = 3'h1 == _T_1246 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2232.6]
  assign _GEN_92 = 3'h2 == _T_1246 ? io_bbLoadOffsets_2 : _GEN_91; // @[LoadQueue.scala 77:20:@2232.6]
  assign _GEN_93 = 3'h3 == _T_1246 ? io_bbLoadOffsets_3 : _GEN_92; // @[LoadQueue.scala 77:20:@2232.6]
  assign _GEN_94 = 3'h4 == _T_1246 ? io_bbLoadOffsets_4 : _GEN_93; // @[LoadQueue.scala 77:20:@2232.6]
  assign _GEN_95 = 3'h5 == _T_1246 ? io_bbLoadOffsets_5 : _GEN_94; // @[LoadQueue.scala 77:20:@2232.6]
  assign _GEN_96 = 3'h6 == _T_1246 ? io_bbLoadOffsets_6 : _GEN_95; // @[LoadQueue.scala 77:20:@2232.6]
  assign _GEN_97 = 3'h7 == _T_1246 ? io_bbLoadOffsets_7 : _GEN_96; // @[LoadQueue.scala 77:20:@2232.6]
  assign _GEN_99 = 3'h1 == _T_1246 ? io_bbLoadPorts_1 : io_bbLoadPorts_0; // @[LoadQueue.scala 78:18:@2239.6]
  assign _GEN_100 = 3'h2 == _T_1246 ? io_bbLoadPorts_2 : _GEN_99; // @[LoadQueue.scala 78:18:@2239.6]
  assign _GEN_101 = 3'h3 == _T_1246 ? 3'h0 : _GEN_100; // @[LoadQueue.scala 78:18:@2239.6]
  assign _GEN_102 = 3'h4 == _T_1246 ? 3'h0 : _GEN_101; // @[LoadQueue.scala 78:18:@2239.6]
  assign _GEN_103 = 3'h5 == _T_1246 ? 3'h0 : _GEN_102; // @[LoadQueue.scala 78:18:@2239.6]
  assign _GEN_104 = 3'h6 == _T_1246 ? 3'h0 : _GEN_103; // @[LoadQueue.scala 78:18:@2239.6]
  assign _GEN_105 = 3'h7 == _T_1246 ? 3'h0 : _GEN_104; // @[LoadQueue.scala 78:18:@2239.6]
  assign _GEN_106 = initBits_5 ? _GEN_97 : offsetQ_5; // @[LoadQueue.scala 76:25:@2225.4]
  assign _GEN_107 = initBits_5 ? _GEN_105 : portQ_5; // @[LoadQueue.scala 76:25:@2225.4]
  assign _T_1264 = _T_1101[2:0]; // @[:@2247.6]
  assign _GEN_109 = 3'h1 == _T_1264 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2248.6]
  assign _GEN_110 = 3'h2 == _T_1264 ? io_bbLoadOffsets_2 : _GEN_109; // @[LoadQueue.scala 77:20:@2248.6]
  assign _GEN_111 = 3'h3 == _T_1264 ? io_bbLoadOffsets_3 : _GEN_110; // @[LoadQueue.scala 77:20:@2248.6]
  assign _GEN_112 = 3'h4 == _T_1264 ? io_bbLoadOffsets_4 : _GEN_111; // @[LoadQueue.scala 77:20:@2248.6]
  assign _GEN_113 = 3'h5 == _T_1264 ? io_bbLoadOffsets_5 : _GEN_112; // @[LoadQueue.scala 77:20:@2248.6]
  assign _GEN_114 = 3'h6 == _T_1264 ? io_bbLoadOffsets_6 : _GEN_113; // @[LoadQueue.scala 77:20:@2248.6]
  assign _GEN_115 = 3'h7 == _T_1264 ? io_bbLoadOffsets_7 : _GEN_114; // @[LoadQueue.scala 77:20:@2248.6]
  assign _GEN_117 = 3'h1 == _T_1264 ? io_bbLoadPorts_1 : io_bbLoadPorts_0; // @[LoadQueue.scala 78:18:@2255.6]
  assign _GEN_118 = 3'h2 == _T_1264 ? io_bbLoadPorts_2 : _GEN_117; // @[LoadQueue.scala 78:18:@2255.6]
  assign _GEN_119 = 3'h3 == _T_1264 ? 3'h0 : _GEN_118; // @[LoadQueue.scala 78:18:@2255.6]
  assign _GEN_120 = 3'h4 == _T_1264 ? 3'h0 : _GEN_119; // @[LoadQueue.scala 78:18:@2255.6]
  assign _GEN_121 = 3'h5 == _T_1264 ? 3'h0 : _GEN_120; // @[LoadQueue.scala 78:18:@2255.6]
  assign _GEN_122 = 3'h6 == _T_1264 ? 3'h0 : _GEN_121; // @[LoadQueue.scala 78:18:@2255.6]
  assign _GEN_123 = 3'h7 == _T_1264 ? 3'h0 : _GEN_122; // @[LoadQueue.scala 78:18:@2255.6]
  assign _GEN_124 = initBits_6 ? _GEN_115 : offsetQ_6; // @[LoadQueue.scala 76:25:@2241.4]
  assign _GEN_125 = initBits_6 ? _GEN_123 : portQ_6; // @[LoadQueue.scala 76:25:@2241.4]
  assign _T_1282 = _T_1110[2:0]; // @[:@2263.6]
  assign _GEN_127 = 3'h1 == _T_1282 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2264.6]
  assign _GEN_128 = 3'h2 == _T_1282 ? io_bbLoadOffsets_2 : _GEN_127; // @[LoadQueue.scala 77:20:@2264.6]
  assign _GEN_129 = 3'h3 == _T_1282 ? io_bbLoadOffsets_3 : _GEN_128; // @[LoadQueue.scala 77:20:@2264.6]
  assign _GEN_130 = 3'h4 == _T_1282 ? io_bbLoadOffsets_4 : _GEN_129; // @[LoadQueue.scala 77:20:@2264.6]
  assign _GEN_131 = 3'h5 == _T_1282 ? io_bbLoadOffsets_5 : _GEN_130; // @[LoadQueue.scala 77:20:@2264.6]
  assign _GEN_132 = 3'h6 == _T_1282 ? io_bbLoadOffsets_6 : _GEN_131; // @[LoadQueue.scala 77:20:@2264.6]
  assign _GEN_133 = 3'h7 == _T_1282 ? io_bbLoadOffsets_7 : _GEN_132; // @[LoadQueue.scala 77:20:@2264.6]
  assign _GEN_135 = 3'h1 == _T_1282 ? io_bbLoadPorts_1 : io_bbLoadPorts_0; // @[LoadQueue.scala 78:18:@2271.6]
  assign _GEN_136 = 3'h2 == _T_1282 ? io_bbLoadPorts_2 : _GEN_135; // @[LoadQueue.scala 78:18:@2271.6]
  assign _GEN_137 = 3'h3 == _T_1282 ? 3'h0 : _GEN_136; // @[LoadQueue.scala 78:18:@2271.6]
  assign _GEN_138 = 3'h4 == _T_1282 ? 3'h0 : _GEN_137; // @[LoadQueue.scala 78:18:@2271.6]
  assign _GEN_139 = 3'h5 == _T_1282 ? 3'h0 : _GEN_138; // @[LoadQueue.scala 78:18:@2271.6]
  assign _GEN_140 = 3'h6 == _T_1282 ? 3'h0 : _GEN_139; // @[LoadQueue.scala 78:18:@2271.6]
  assign _GEN_141 = 3'h7 == _T_1282 ? 3'h0 : _GEN_140; // @[LoadQueue.scala 78:18:@2271.6]
  assign _GEN_142 = initBits_7 ? _GEN_133 : offsetQ_7; // @[LoadQueue.scala 76:25:@2257.4]
  assign _GEN_143 = initBits_7 ? _GEN_141 : portQ_7; // @[LoadQueue.scala 76:25:@2257.4]
  assign _T_1304 = _GEN_7 + 3'h1; // @[util.scala 10:8:@2282.6]
  assign _GEN_72 = _T_1304 % 4'h8; // @[util.scala 10:14:@2283.6]
  assign _T_1305 = _GEN_72[3:0]; // @[util.scala 10:14:@2283.6]
  assign _GEN_799 = {{1'd0}, io_storeTail}; // @[LoadQueue.scala 97:56:@2284.6]
  assign _T_1306 = _T_1305 == _GEN_799; // @[LoadQueue.scala 97:56:@2284.6]
  assign _T_1307 = io_storeEmpty & _T_1306; // @[LoadQueue.scala 96:50:@2285.6]
  assign _T_1309 = _T_1307 == 1'h0; // @[LoadQueue.scala 96:34:@2286.6]
  assign _T_1311 = previousStoreHead <= offsetQ_0; // @[LoadQueue.scala 101:36:@2294.8]
  assign _T_1312 = offsetQ_0 < io_storeHead; // @[LoadQueue.scala 101:86:@2295.8]
  assign _T_1313 = _T_1311 & _T_1312; // @[LoadQueue.scala 101:61:@2296.8]
  assign _T_1315 = previousStoreHead > io_storeHead; // @[LoadQueue.scala 103:36:@2301.10]
  assign _T_1316 = io_storeHead <= offsetQ_0; // @[LoadQueue.scala 103:69:@2302.10]
  assign _T_1317 = offsetQ_0 < previousStoreHead; // @[LoadQueue.scala 104:31:@2303.10]
  assign _T_1318 = _T_1316 & _T_1317; // @[LoadQueue.scala 103:94:@2304.10]
  assign _T_1320 = _T_1318 == 1'h0; // @[LoadQueue.scala 103:54:@2305.10]
  assign _T_1321 = _T_1315 & _T_1320; // @[LoadQueue.scala 103:51:@2306.10]
  assign _GEN_152 = _T_1321 ? 1'h0 : checkBits_0; // @[LoadQueue.scala 104:53:@2307.10]
  assign _GEN_153 = _T_1313 ? 1'h0 : _GEN_152; // @[LoadQueue.scala 101:102:@2297.8]
  assign _GEN_154 = io_storeEmpty ? 1'h0 : _GEN_153; // @[LoadQueue.scala 99:27:@2290.6]
  assign _GEN_155 = initBits_0 ? _T_1309 : _GEN_154; // @[LoadQueue.scala 95:34:@2275.4]
  assign _T_1334 = _GEN_25 + 3'h1; // @[util.scala 10:8:@2318.6]
  assign _GEN_80 = _T_1334 % 4'h8; // @[util.scala 10:14:@2319.6]
  assign _T_1335 = _GEN_80[3:0]; // @[util.scala 10:14:@2319.6]
  assign _T_1336 = _T_1335 == _GEN_799; // @[LoadQueue.scala 97:56:@2320.6]
  assign _T_1337 = io_storeEmpty & _T_1336; // @[LoadQueue.scala 96:50:@2321.6]
  assign _T_1339 = _T_1337 == 1'h0; // @[LoadQueue.scala 96:34:@2322.6]
  assign _T_1341 = previousStoreHead <= offsetQ_1; // @[LoadQueue.scala 101:36:@2330.8]
  assign _T_1342 = offsetQ_1 < io_storeHead; // @[LoadQueue.scala 101:86:@2331.8]
  assign _T_1343 = _T_1341 & _T_1342; // @[LoadQueue.scala 101:61:@2332.8]
  assign _T_1346 = io_storeHead <= offsetQ_1; // @[LoadQueue.scala 103:69:@2338.10]
  assign _T_1347 = offsetQ_1 < previousStoreHead; // @[LoadQueue.scala 104:31:@2339.10]
  assign _T_1348 = _T_1346 & _T_1347; // @[LoadQueue.scala 103:94:@2340.10]
  assign _T_1350 = _T_1348 == 1'h0; // @[LoadQueue.scala 103:54:@2341.10]
  assign _T_1351 = _T_1315 & _T_1350; // @[LoadQueue.scala 103:51:@2342.10]
  assign _GEN_164 = _T_1351 ? 1'h0 : checkBits_1; // @[LoadQueue.scala 104:53:@2343.10]
  assign _GEN_165 = _T_1343 ? 1'h0 : _GEN_164; // @[LoadQueue.scala 101:102:@2333.8]
  assign _GEN_166 = io_storeEmpty ? 1'h0 : _GEN_165; // @[LoadQueue.scala 99:27:@2326.6]
  assign _GEN_167 = initBits_1 ? _T_1339 : _GEN_166; // @[LoadQueue.scala 95:34:@2311.4]
  assign _T_1364 = _GEN_43 + 3'h1; // @[util.scala 10:8:@2354.6]
  assign _GEN_90 = _T_1364 % 4'h8; // @[util.scala 10:14:@2355.6]
  assign _T_1365 = _GEN_90[3:0]; // @[util.scala 10:14:@2355.6]
  assign _T_1366 = _T_1365 == _GEN_799; // @[LoadQueue.scala 97:56:@2356.6]
  assign _T_1367 = io_storeEmpty & _T_1366; // @[LoadQueue.scala 96:50:@2357.6]
  assign _T_1369 = _T_1367 == 1'h0; // @[LoadQueue.scala 96:34:@2358.6]
  assign _T_1371 = previousStoreHead <= offsetQ_2; // @[LoadQueue.scala 101:36:@2366.8]
  assign _T_1372 = offsetQ_2 < io_storeHead; // @[LoadQueue.scala 101:86:@2367.8]
  assign _T_1373 = _T_1371 & _T_1372; // @[LoadQueue.scala 101:61:@2368.8]
  assign _T_1376 = io_storeHead <= offsetQ_2; // @[LoadQueue.scala 103:69:@2374.10]
  assign _T_1377 = offsetQ_2 < previousStoreHead; // @[LoadQueue.scala 104:31:@2375.10]
  assign _T_1378 = _T_1376 & _T_1377; // @[LoadQueue.scala 103:94:@2376.10]
  assign _T_1380 = _T_1378 == 1'h0; // @[LoadQueue.scala 103:54:@2377.10]
  assign _T_1381 = _T_1315 & _T_1380; // @[LoadQueue.scala 103:51:@2378.10]
  assign _GEN_176 = _T_1381 ? 1'h0 : checkBits_2; // @[LoadQueue.scala 104:53:@2379.10]
  assign _GEN_177 = _T_1373 ? 1'h0 : _GEN_176; // @[LoadQueue.scala 101:102:@2369.8]
  assign _GEN_178 = io_storeEmpty ? 1'h0 : _GEN_177; // @[LoadQueue.scala 99:27:@2362.6]
  assign _GEN_179 = initBits_2 ? _T_1369 : _GEN_178; // @[LoadQueue.scala 95:34:@2347.4]
  assign _T_1394 = _GEN_61 + 3'h1; // @[util.scala 10:8:@2390.6]
  assign _GEN_98 = _T_1394 % 4'h8; // @[util.scala 10:14:@2391.6]
  assign _T_1395 = _GEN_98[3:0]; // @[util.scala 10:14:@2391.6]
  assign _T_1396 = _T_1395 == _GEN_799; // @[LoadQueue.scala 97:56:@2392.6]
  assign _T_1397 = io_storeEmpty & _T_1396; // @[LoadQueue.scala 96:50:@2393.6]
  assign _T_1399 = _T_1397 == 1'h0; // @[LoadQueue.scala 96:34:@2394.6]
  assign _T_1401 = previousStoreHead <= offsetQ_3; // @[LoadQueue.scala 101:36:@2402.8]
  assign _T_1402 = offsetQ_3 < io_storeHead; // @[LoadQueue.scala 101:86:@2403.8]
  assign _T_1403 = _T_1401 & _T_1402; // @[LoadQueue.scala 101:61:@2404.8]
  assign _T_1406 = io_storeHead <= offsetQ_3; // @[LoadQueue.scala 103:69:@2410.10]
  assign _T_1407 = offsetQ_3 < previousStoreHead; // @[LoadQueue.scala 104:31:@2411.10]
  assign _T_1408 = _T_1406 & _T_1407; // @[LoadQueue.scala 103:94:@2412.10]
  assign _T_1410 = _T_1408 == 1'h0; // @[LoadQueue.scala 103:54:@2413.10]
  assign _T_1411 = _T_1315 & _T_1410; // @[LoadQueue.scala 103:51:@2414.10]
  assign _GEN_188 = _T_1411 ? 1'h0 : checkBits_3; // @[LoadQueue.scala 104:53:@2415.10]
  assign _GEN_189 = _T_1403 ? 1'h0 : _GEN_188; // @[LoadQueue.scala 101:102:@2405.8]
  assign _GEN_190 = io_storeEmpty ? 1'h0 : _GEN_189; // @[LoadQueue.scala 99:27:@2398.6]
  assign _GEN_191 = initBits_3 ? _T_1399 : _GEN_190; // @[LoadQueue.scala 95:34:@2383.4]
  assign _T_1424 = _GEN_79 + 3'h1; // @[util.scala 10:8:@2426.6]
  assign _GEN_108 = _T_1424 % 4'h8; // @[util.scala 10:14:@2427.6]
  assign _T_1425 = _GEN_108[3:0]; // @[util.scala 10:14:@2427.6]
  assign _T_1426 = _T_1425 == _GEN_799; // @[LoadQueue.scala 97:56:@2428.6]
  assign _T_1427 = io_storeEmpty & _T_1426; // @[LoadQueue.scala 96:50:@2429.6]
  assign _T_1429 = _T_1427 == 1'h0; // @[LoadQueue.scala 96:34:@2430.6]
  assign _T_1431 = previousStoreHead <= offsetQ_4; // @[LoadQueue.scala 101:36:@2438.8]
  assign _T_1432 = offsetQ_4 < io_storeHead; // @[LoadQueue.scala 101:86:@2439.8]
  assign _T_1433 = _T_1431 & _T_1432; // @[LoadQueue.scala 101:61:@2440.8]
  assign _T_1436 = io_storeHead <= offsetQ_4; // @[LoadQueue.scala 103:69:@2446.10]
  assign _T_1437 = offsetQ_4 < previousStoreHead; // @[LoadQueue.scala 104:31:@2447.10]
  assign _T_1438 = _T_1436 & _T_1437; // @[LoadQueue.scala 103:94:@2448.10]
  assign _T_1440 = _T_1438 == 1'h0; // @[LoadQueue.scala 103:54:@2449.10]
  assign _T_1441 = _T_1315 & _T_1440; // @[LoadQueue.scala 103:51:@2450.10]
  assign _GEN_200 = _T_1441 ? 1'h0 : checkBits_4; // @[LoadQueue.scala 104:53:@2451.10]
  assign _GEN_201 = _T_1433 ? 1'h0 : _GEN_200; // @[LoadQueue.scala 101:102:@2441.8]
  assign _GEN_202 = io_storeEmpty ? 1'h0 : _GEN_201; // @[LoadQueue.scala 99:27:@2434.6]
  assign _GEN_203 = initBits_4 ? _T_1429 : _GEN_202; // @[LoadQueue.scala 95:34:@2419.4]
  assign _T_1454 = _GEN_97 + 3'h1; // @[util.scala 10:8:@2462.6]
  assign _GEN_116 = _T_1454 % 4'h8; // @[util.scala 10:14:@2463.6]
  assign _T_1455 = _GEN_116[3:0]; // @[util.scala 10:14:@2463.6]
  assign _T_1456 = _T_1455 == _GEN_799; // @[LoadQueue.scala 97:56:@2464.6]
  assign _T_1457 = io_storeEmpty & _T_1456; // @[LoadQueue.scala 96:50:@2465.6]
  assign _T_1459 = _T_1457 == 1'h0; // @[LoadQueue.scala 96:34:@2466.6]
  assign _T_1461 = previousStoreHead <= offsetQ_5; // @[LoadQueue.scala 101:36:@2474.8]
  assign _T_1462 = offsetQ_5 < io_storeHead; // @[LoadQueue.scala 101:86:@2475.8]
  assign _T_1463 = _T_1461 & _T_1462; // @[LoadQueue.scala 101:61:@2476.8]
  assign _T_1466 = io_storeHead <= offsetQ_5; // @[LoadQueue.scala 103:69:@2482.10]
  assign _T_1467 = offsetQ_5 < previousStoreHead; // @[LoadQueue.scala 104:31:@2483.10]
  assign _T_1468 = _T_1466 & _T_1467; // @[LoadQueue.scala 103:94:@2484.10]
  assign _T_1470 = _T_1468 == 1'h0; // @[LoadQueue.scala 103:54:@2485.10]
  assign _T_1471 = _T_1315 & _T_1470; // @[LoadQueue.scala 103:51:@2486.10]
  assign _GEN_212 = _T_1471 ? 1'h0 : checkBits_5; // @[LoadQueue.scala 104:53:@2487.10]
  assign _GEN_213 = _T_1463 ? 1'h0 : _GEN_212; // @[LoadQueue.scala 101:102:@2477.8]
  assign _GEN_214 = io_storeEmpty ? 1'h0 : _GEN_213; // @[LoadQueue.scala 99:27:@2470.6]
  assign _GEN_215 = initBits_5 ? _T_1459 : _GEN_214; // @[LoadQueue.scala 95:34:@2455.4]
  assign _T_1484 = _GEN_115 + 3'h1; // @[util.scala 10:8:@2498.6]
  assign _GEN_126 = _T_1484 % 4'h8; // @[util.scala 10:14:@2499.6]
  assign _T_1485 = _GEN_126[3:0]; // @[util.scala 10:14:@2499.6]
  assign _T_1486 = _T_1485 == _GEN_799; // @[LoadQueue.scala 97:56:@2500.6]
  assign _T_1487 = io_storeEmpty & _T_1486; // @[LoadQueue.scala 96:50:@2501.6]
  assign _T_1489 = _T_1487 == 1'h0; // @[LoadQueue.scala 96:34:@2502.6]
  assign _T_1491 = previousStoreHead <= offsetQ_6; // @[LoadQueue.scala 101:36:@2510.8]
  assign _T_1492 = offsetQ_6 < io_storeHead; // @[LoadQueue.scala 101:86:@2511.8]
  assign _T_1493 = _T_1491 & _T_1492; // @[LoadQueue.scala 101:61:@2512.8]
  assign _T_1496 = io_storeHead <= offsetQ_6; // @[LoadQueue.scala 103:69:@2518.10]
  assign _T_1497 = offsetQ_6 < previousStoreHead; // @[LoadQueue.scala 104:31:@2519.10]
  assign _T_1498 = _T_1496 & _T_1497; // @[LoadQueue.scala 103:94:@2520.10]
  assign _T_1500 = _T_1498 == 1'h0; // @[LoadQueue.scala 103:54:@2521.10]
  assign _T_1501 = _T_1315 & _T_1500; // @[LoadQueue.scala 103:51:@2522.10]
  assign _GEN_224 = _T_1501 ? 1'h0 : checkBits_6; // @[LoadQueue.scala 104:53:@2523.10]
  assign _GEN_225 = _T_1493 ? 1'h0 : _GEN_224; // @[LoadQueue.scala 101:102:@2513.8]
  assign _GEN_226 = io_storeEmpty ? 1'h0 : _GEN_225; // @[LoadQueue.scala 99:27:@2506.6]
  assign _GEN_227 = initBits_6 ? _T_1489 : _GEN_226; // @[LoadQueue.scala 95:34:@2491.4]
  assign _T_1514 = _GEN_133 + 3'h1; // @[util.scala 10:8:@2534.6]
  assign _GEN_134 = _T_1514 % 4'h8; // @[util.scala 10:14:@2535.6]
  assign _T_1515 = _GEN_134[3:0]; // @[util.scala 10:14:@2535.6]
  assign _T_1516 = _T_1515 == _GEN_799; // @[LoadQueue.scala 97:56:@2536.6]
  assign _T_1517 = io_storeEmpty & _T_1516; // @[LoadQueue.scala 96:50:@2537.6]
  assign _T_1519 = _T_1517 == 1'h0; // @[LoadQueue.scala 96:34:@2538.6]
  assign _T_1521 = previousStoreHead <= offsetQ_7; // @[LoadQueue.scala 101:36:@2546.8]
  assign _T_1522 = offsetQ_7 < io_storeHead; // @[LoadQueue.scala 101:86:@2547.8]
  assign _T_1523 = _T_1521 & _T_1522; // @[LoadQueue.scala 101:61:@2548.8]
  assign _T_1526 = io_storeHead <= offsetQ_7; // @[LoadQueue.scala 103:69:@2554.10]
  assign _T_1527 = offsetQ_7 < previousStoreHead; // @[LoadQueue.scala 104:31:@2555.10]
  assign _T_1528 = _T_1526 & _T_1527; // @[LoadQueue.scala 103:94:@2556.10]
  assign _T_1530 = _T_1528 == 1'h0; // @[LoadQueue.scala 103:54:@2557.10]
  assign _T_1531 = _T_1315 & _T_1530; // @[LoadQueue.scala 103:51:@2558.10]
  assign _GEN_236 = _T_1531 ? 1'h0 : checkBits_7; // @[LoadQueue.scala 104:53:@2559.10]
  assign _GEN_237 = _T_1523 ? 1'h0 : _GEN_236; // @[LoadQueue.scala 101:102:@2549.8]
  assign _GEN_238 = io_storeEmpty ? 1'h0 : _GEN_237; // @[LoadQueue.scala 99:27:@2542.6]
  assign _GEN_239 = initBits_7 ? _T_1519 : _GEN_238; // @[LoadQueue.scala 95:34:@2527.4]
  assign _T_1535 = 8'h1 << io_storeHead; // @[OneHot.scala 52:12:@2564.4]
  assign _T_1537 = _T_1535[0]; // @[util.scala 60:60:@2566.4]
  assign _T_1538 = _T_1535[1]; // @[util.scala 60:60:@2567.4]
  assign _T_1539 = _T_1535[2]; // @[util.scala 60:60:@2568.4]
  assign _T_1540 = _T_1535[3]; // @[util.scala 60:60:@2569.4]
  assign _T_1541 = _T_1535[4]; // @[util.scala 60:60:@2570.4]
  assign _T_1542 = _T_1535[5]; // @[util.scala 60:60:@2571.4]
  assign _T_1543 = _T_1535[6]; // @[util.scala 60:60:@2572.4]
  assign _T_1544 = _T_1535[7]; // @[util.scala 60:60:@2573.4]
  assign _T_2323 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0}; // @[Mux.scala 19:72:@3025.4]
  assign _T_2325 = _T_1537 ? _T_2323 : 256'h0; // @[Mux.scala 19:72:@3026.4]
  assign _T_2332 = {io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1}; // @[Mux.scala 19:72:@3033.4]
  assign _T_2334 = _T_1538 ? _T_2332 : 256'h0; // @[Mux.scala 19:72:@3034.4]
  assign _T_2341 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2}; // @[Mux.scala 19:72:@3041.4]
  assign _T_2343 = _T_1539 ? _T_2341 : 256'h0; // @[Mux.scala 19:72:@3042.4]
  assign _T_2350 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3}; // @[Mux.scala 19:72:@3049.4]
  assign _T_2352 = _T_1540 ? _T_2350 : 256'h0; // @[Mux.scala 19:72:@3050.4]
  assign _T_2359 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4}; // @[Mux.scala 19:72:@3057.4]
  assign _T_2361 = _T_1541 ? _T_2359 : 256'h0; // @[Mux.scala 19:72:@3058.4]
  assign _T_2368 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5}; // @[Mux.scala 19:72:@3065.4]
  assign _T_2370 = _T_1542 ? _T_2368 : 256'h0; // @[Mux.scala 19:72:@3066.4]
  assign _T_2377 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6}; // @[Mux.scala 19:72:@3073.4]
  assign _T_2379 = _T_1543 ? _T_2377 : 256'h0; // @[Mux.scala 19:72:@3074.4]
  assign _T_2386 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7}; // @[Mux.scala 19:72:@3081.4]
  assign _T_2388 = _T_1544 ? _T_2386 : 256'h0; // @[Mux.scala 19:72:@3082.4]
  assign _T_2389 = _T_2325 | _T_2334; // @[Mux.scala 19:72:@3083.4]
  assign _T_2390 = _T_2389 | _T_2343; // @[Mux.scala 19:72:@3084.4]
  assign _T_2391 = _T_2390 | _T_2352; // @[Mux.scala 19:72:@3085.4]
  assign _T_2392 = _T_2391 | _T_2361; // @[Mux.scala 19:72:@3086.4]
  assign _T_2393 = _T_2392 | _T_2370; // @[Mux.scala 19:72:@3087.4]
  assign _T_2394 = _T_2393 | _T_2379; // @[Mux.scala 19:72:@3088.4]
  assign _T_2395 = _T_2394 | _T_2388; // @[Mux.scala 19:72:@3089.4]
  assign _T_2636 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0}; // @[Mux.scala 19:72:@3207.4]
  assign _T_2638 = _T_1537 ? _T_2636 : 8'h0; // @[Mux.scala 19:72:@3208.4]
  assign _T_2645 = {io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1}; // @[Mux.scala 19:72:@3215.4]
  assign _T_2647 = _T_1538 ? _T_2645 : 8'h0; // @[Mux.scala 19:72:@3216.4]
  assign _T_2654 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2}; // @[Mux.scala 19:72:@3223.4]
  assign _T_2656 = _T_1539 ? _T_2654 : 8'h0; // @[Mux.scala 19:72:@3224.4]
  assign _T_2663 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3}; // @[Mux.scala 19:72:@3231.4]
  assign _T_2665 = _T_1540 ? _T_2663 : 8'h0; // @[Mux.scala 19:72:@3232.4]
  assign _T_2672 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4}; // @[Mux.scala 19:72:@3239.4]
  assign _T_2674 = _T_1541 ? _T_2672 : 8'h0; // @[Mux.scala 19:72:@3240.4]
  assign _T_2681 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5}; // @[Mux.scala 19:72:@3247.4]
  assign _T_2683 = _T_1542 ? _T_2681 : 8'h0; // @[Mux.scala 19:72:@3248.4]
  assign _T_2690 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6}; // @[Mux.scala 19:72:@3255.4]
  assign _T_2692 = _T_1543 ? _T_2690 : 8'h0; // @[Mux.scala 19:72:@3256.4]
  assign _T_2699 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7}; // @[Mux.scala 19:72:@3263.4]
  assign _T_2701 = _T_1544 ? _T_2699 : 8'h0; // @[Mux.scala 19:72:@3264.4]
  assign _T_2702 = _T_2638 | _T_2647; // @[Mux.scala 19:72:@3265.4]
  assign _T_2703 = _T_2702 | _T_2656; // @[Mux.scala 19:72:@3266.4]
  assign _T_2704 = _T_2703 | _T_2665; // @[Mux.scala 19:72:@3267.4]
  assign _T_2705 = _T_2704 | _T_2674; // @[Mux.scala 19:72:@3268.4]
  assign _T_2706 = _T_2705 | _T_2683; // @[Mux.scala 19:72:@3269.4]
  assign _T_2707 = _T_2706 | _T_2692; // @[Mux.scala 19:72:@3270.4]
  assign _T_2708 = _T_2707 | _T_2701; // @[Mux.scala 19:72:@3271.4]
  assign _T_2785 = io_storeHead < io_storeTail; // @[LoadQueue.scala 121:105:@3291.4]
  assign _T_2787 = io_storeHead <= 3'h0; // @[LoadQueue.scala 122:18:@3292.4]
  assign _T_2789 = 3'h0 < io_storeTail; // @[LoadQueue.scala 122:36:@3293.4]
  assign _T_2790 = _T_2787 & _T_2789; // @[LoadQueue.scala 122:27:@3294.4]
  assign _T_2792 = io_storeEmpty == 1'h0; // @[LoadQueue.scala 122:52:@3295.4]
  assign _T_2794 = io_storeTail <= 3'h0; // @[LoadQueue.scala 122:85:@3296.4]
  assign _T_2796 = 3'h0 < io_storeHead; // @[LoadQueue.scala 122:103:@3297.4]
  assign _T_2797 = _T_2794 & _T_2796; // @[LoadQueue.scala 122:94:@3298.4]
  assign _T_2799 = _T_2797 == 1'h0; // @[LoadQueue.scala 122:70:@3299.4]
  assign _T_2800 = _T_2792 & _T_2799; // @[LoadQueue.scala 122:67:@3300.4]
  assign validEntriesInStoreQ_0 = _T_2785 ? _T_2790 : _T_2800; // @[LoadQueue.scala 121:91:@3301.4]
  assign _T_2804 = io_storeHead <= 3'h1; // @[LoadQueue.scala 122:18:@3303.4]
  assign _T_2806 = 3'h1 < io_storeTail; // @[LoadQueue.scala 122:36:@3304.4]
  assign _T_2807 = _T_2804 & _T_2806; // @[LoadQueue.scala 122:27:@3305.4]
  assign _T_2811 = io_storeTail <= 3'h1; // @[LoadQueue.scala 122:85:@3307.4]
  assign _T_2813 = 3'h1 < io_storeHead; // @[LoadQueue.scala 122:103:@3308.4]
  assign _T_2814 = _T_2811 & _T_2813; // @[LoadQueue.scala 122:94:@3309.4]
  assign _T_2816 = _T_2814 == 1'h0; // @[LoadQueue.scala 122:70:@3310.4]
  assign _T_2817 = _T_2792 & _T_2816; // @[LoadQueue.scala 122:67:@3311.4]
  assign validEntriesInStoreQ_1 = _T_2785 ? _T_2807 : _T_2817; // @[LoadQueue.scala 121:91:@3312.4]
  assign _T_2821 = io_storeHead <= 3'h2; // @[LoadQueue.scala 122:18:@3314.4]
  assign _T_2823 = 3'h2 < io_storeTail; // @[LoadQueue.scala 122:36:@3315.4]
  assign _T_2824 = _T_2821 & _T_2823; // @[LoadQueue.scala 122:27:@3316.4]
  assign _T_2828 = io_storeTail <= 3'h2; // @[LoadQueue.scala 122:85:@3318.4]
  assign _T_2830 = 3'h2 < io_storeHead; // @[LoadQueue.scala 122:103:@3319.4]
  assign _T_2831 = _T_2828 & _T_2830; // @[LoadQueue.scala 122:94:@3320.4]
  assign _T_2833 = _T_2831 == 1'h0; // @[LoadQueue.scala 122:70:@3321.4]
  assign _T_2834 = _T_2792 & _T_2833; // @[LoadQueue.scala 122:67:@3322.4]
  assign validEntriesInStoreQ_2 = _T_2785 ? _T_2824 : _T_2834; // @[LoadQueue.scala 121:91:@3323.4]
  assign _T_2838 = io_storeHead <= 3'h3; // @[LoadQueue.scala 122:18:@3325.4]
  assign _T_2840 = 3'h3 < io_storeTail; // @[LoadQueue.scala 122:36:@3326.4]
  assign _T_2841 = _T_2838 & _T_2840; // @[LoadQueue.scala 122:27:@3327.4]
  assign _T_2845 = io_storeTail <= 3'h3; // @[LoadQueue.scala 122:85:@3329.4]
  assign _T_2847 = 3'h3 < io_storeHead; // @[LoadQueue.scala 122:103:@3330.4]
  assign _T_2848 = _T_2845 & _T_2847; // @[LoadQueue.scala 122:94:@3331.4]
  assign _T_2850 = _T_2848 == 1'h0; // @[LoadQueue.scala 122:70:@3332.4]
  assign _T_2851 = _T_2792 & _T_2850; // @[LoadQueue.scala 122:67:@3333.4]
  assign validEntriesInStoreQ_3 = _T_2785 ? _T_2841 : _T_2851; // @[LoadQueue.scala 121:91:@3334.4]
  assign _T_2855 = io_storeHead <= 3'h4; // @[LoadQueue.scala 122:18:@3336.4]
  assign _T_2857 = 3'h4 < io_storeTail; // @[LoadQueue.scala 122:36:@3337.4]
  assign _T_2858 = _T_2855 & _T_2857; // @[LoadQueue.scala 122:27:@3338.4]
  assign _T_2862 = io_storeTail <= 3'h4; // @[LoadQueue.scala 122:85:@3340.4]
  assign _T_2864 = 3'h4 < io_storeHead; // @[LoadQueue.scala 122:103:@3341.4]
  assign _T_2865 = _T_2862 & _T_2864; // @[LoadQueue.scala 122:94:@3342.4]
  assign _T_2867 = _T_2865 == 1'h0; // @[LoadQueue.scala 122:70:@3343.4]
  assign _T_2868 = _T_2792 & _T_2867; // @[LoadQueue.scala 122:67:@3344.4]
  assign validEntriesInStoreQ_4 = _T_2785 ? _T_2858 : _T_2868; // @[LoadQueue.scala 121:91:@3345.4]
  assign _T_2872 = io_storeHead <= 3'h5; // @[LoadQueue.scala 122:18:@3347.4]
  assign _T_2874 = 3'h5 < io_storeTail; // @[LoadQueue.scala 122:36:@3348.4]
  assign _T_2875 = _T_2872 & _T_2874; // @[LoadQueue.scala 122:27:@3349.4]
  assign _T_2879 = io_storeTail <= 3'h5; // @[LoadQueue.scala 122:85:@3351.4]
  assign _T_2881 = 3'h5 < io_storeHead; // @[LoadQueue.scala 122:103:@3352.4]
  assign _T_2882 = _T_2879 & _T_2881; // @[LoadQueue.scala 122:94:@3353.4]
  assign _T_2884 = _T_2882 == 1'h0; // @[LoadQueue.scala 122:70:@3354.4]
  assign _T_2885 = _T_2792 & _T_2884; // @[LoadQueue.scala 122:67:@3355.4]
  assign validEntriesInStoreQ_5 = _T_2785 ? _T_2875 : _T_2885; // @[LoadQueue.scala 121:91:@3356.4]
  assign _T_2889 = io_storeHead <= 3'h6; // @[LoadQueue.scala 122:18:@3358.4]
  assign _T_2891 = 3'h6 < io_storeTail; // @[LoadQueue.scala 122:36:@3359.4]
  assign _T_2892 = _T_2889 & _T_2891; // @[LoadQueue.scala 122:27:@3360.4]
  assign _T_2896 = io_storeTail <= 3'h6; // @[LoadQueue.scala 122:85:@3362.4]
  assign _T_2898 = 3'h6 < io_storeHead; // @[LoadQueue.scala 122:103:@3363.4]
  assign _T_2899 = _T_2896 & _T_2898; // @[LoadQueue.scala 122:94:@3364.4]
  assign _T_2901 = _T_2899 == 1'h0; // @[LoadQueue.scala 122:70:@3365.4]
  assign _T_2902 = _T_2792 & _T_2901; // @[LoadQueue.scala 122:67:@3366.4]
  assign validEntriesInStoreQ_6 = _T_2785 ? _T_2892 : _T_2902; // @[LoadQueue.scala 121:91:@3367.4]
  assign validEntriesInStoreQ_7 = _T_2785 ? 1'h0 : _T_2792; // @[LoadQueue.scala 121:91:@3378.4]
  assign storesToCheck_0_0 = _T_1316 ? _T_2787 : 1'h1; // @[LoadQueue.scala 131:10:@3397.4]
  assign _T_3318 = 3'h1 <= offsetQ_0; // @[LoadQueue.scala 131:81:@3400.4]
  assign _T_3319 = _T_2804 & _T_3318; // @[LoadQueue.scala 131:72:@3401.4]
  assign _T_3321 = offsetQ_0 < 3'h1; // @[LoadQueue.scala 132:33:@3402.4]
  assign _T_3324 = _T_3321 & _T_2813; // @[LoadQueue.scala 132:41:@3404.4]
  assign _T_3326 = _T_3324 == 1'h0; // @[LoadQueue.scala 132:9:@3405.4]
  assign storesToCheck_0_1 = _T_1316 ? _T_3319 : _T_3326; // @[LoadQueue.scala 131:10:@3406.4]
  assign _T_3332 = 3'h2 <= offsetQ_0; // @[LoadQueue.scala 131:81:@3409.4]
  assign _T_3333 = _T_2821 & _T_3332; // @[LoadQueue.scala 131:72:@3410.4]
  assign _T_3335 = offsetQ_0 < 3'h2; // @[LoadQueue.scala 132:33:@3411.4]
  assign _T_3338 = _T_3335 & _T_2830; // @[LoadQueue.scala 132:41:@3413.4]
  assign _T_3340 = _T_3338 == 1'h0; // @[LoadQueue.scala 132:9:@3414.4]
  assign storesToCheck_0_2 = _T_1316 ? _T_3333 : _T_3340; // @[LoadQueue.scala 131:10:@3415.4]
  assign _T_3346 = 3'h3 <= offsetQ_0; // @[LoadQueue.scala 131:81:@3418.4]
  assign _T_3347 = _T_2838 & _T_3346; // @[LoadQueue.scala 131:72:@3419.4]
  assign _T_3349 = offsetQ_0 < 3'h3; // @[LoadQueue.scala 132:33:@3420.4]
  assign _T_3352 = _T_3349 & _T_2847; // @[LoadQueue.scala 132:41:@3422.4]
  assign _T_3354 = _T_3352 == 1'h0; // @[LoadQueue.scala 132:9:@3423.4]
  assign storesToCheck_0_3 = _T_1316 ? _T_3347 : _T_3354; // @[LoadQueue.scala 131:10:@3424.4]
  assign _T_3360 = 3'h4 <= offsetQ_0; // @[LoadQueue.scala 131:81:@3427.4]
  assign _T_3361 = _T_2855 & _T_3360; // @[LoadQueue.scala 131:72:@3428.4]
  assign _T_3363 = offsetQ_0 < 3'h4; // @[LoadQueue.scala 132:33:@3429.4]
  assign _T_3366 = _T_3363 & _T_2864; // @[LoadQueue.scala 132:41:@3431.4]
  assign _T_3368 = _T_3366 == 1'h0; // @[LoadQueue.scala 132:9:@3432.4]
  assign storesToCheck_0_4 = _T_1316 ? _T_3361 : _T_3368; // @[LoadQueue.scala 131:10:@3433.4]
  assign _T_3374 = 3'h5 <= offsetQ_0; // @[LoadQueue.scala 131:81:@3436.4]
  assign _T_3375 = _T_2872 & _T_3374; // @[LoadQueue.scala 131:72:@3437.4]
  assign _T_3377 = offsetQ_0 < 3'h5; // @[LoadQueue.scala 132:33:@3438.4]
  assign _T_3380 = _T_3377 & _T_2881; // @[LoadQueue.scala 132:41:@3440.4]
  assign _T_3382 = _T_3380 == 1'h0; // @[LoadQueue.scala 132:9:@3441.4]
  assign storesToCheck_0_5 = _T_1316 ? _T_3375 : _T_3382; // @[LoadQueue.scala 131:10:@3442.4]
  assign _T_3388 = 3'h6 <= offsetQ_0; // @[LoadQueue.scala 131:81:@3445.4]
  assign _T_3389 = _T_2889 & _T_3388; // @[LoadQueue.scala 131:72:@3446.4]
  assign _T_3391 = offsetQ_0 < 3'h6; // @[LoadQueue.scala 132:33:@3447.4]
  assign _T_3394 = _T_3391 & _T_2898; // @[LoadQueue.scala 132:41:@3449.4]
  assign _T_3396 = _T_3394 == 1'h0; // @[LoadQueue.scala 132:9:@3450.4]
  assign storesToCheck_0_6 = _T_1316 ? _T_3389 : _T_3396; // @[LoadQueue.scala 131:10:@3451.4]
  assign _T_3402 = 3'h7 <= offsetQ_0; // @[LoadQueue.scala 131:81:@3454.4]
  assign storesToCheck_0_7 = _T_1316 ? _T_3402 : 1'h1; // @[LoadQueue.scala 131:10:@3460.4]
  assign storesToCheck_1_0 = _T_1346 ? _T_2787 : 1'h1; // @[LoadQueue.scala 131:10:@3486.4]
  assign _T_3444 = 3'h1 <= offsetQ_1; // @[LoadQueue.scala 131:81:@3489.4]
  assign _T_3445 = _T_2804 & _T_3444; // @[LoadQueue.scala 131:72:@3490.4]
  assign _T_3447 = offsetQ_1 < 3'h1; // @[LoadQueue.scala 132:33:@3491.4]
  assign _T_3450 = _T_3447 & _T_2813; // @[LoadQueue.scala 132:41:@3493.4]
  assign _T_3452 = _T_3450 == 1'h0; // @[LoadQueue.scala 132:9:@3494.4]
  assign storesToCheck_1_1 = _T_1346 ? _T_3445 : _T_3452; // @[LoadQueue.scala 131:10:@3495.4]
  assign _T_3458 = 3'h2 <= offsetQ_1; // @[LoadQueue.scala 131:81:@3498.4]
  assign _T_3459 = _T_2821 & _T_3458; // @[LoadQueue.scala 131:72:@3499.4]
  assign _T_3461 = offsetQ_1 < 3'h2; // @[LoadQueue.scala 132:33:@3500.4]
  assign _T_3464 = _T_3461 & _T_2830; // @[LoadQueue.scala 132:41:@3502.4]
  assign _T_3466 = _T_3464 == 1'h0; // @[LoadQueue.scala 132:9:@3503.4]
  assign storesToCheck_1_2 = _T_1346 ? _T_3459 : _T_3466; // @[LoadQueue.scala 131:10:@3504.4]
  assign _T_3472 = 3'h3 <= offsetQ_1; // @[LoadQueue.scala 131:81:@3507.4]
  assign _T_3473 = _T_2838 & _T_3472; // @[LoadQueue.scala 131:72:@3508.4]
  assign _T_3475 = offsetQ_1 < 3'h3; // @[LoadQueue.scala 132:33:@3509.4]
  assign _T_3478 = _T_3475 & _T_2847; // @[LoadQueue.scala 132:41:@3511.4]
  assign _T_3480 = _T_3478 == 1'h0; // @[LoadQueue.scala 132:9:@3512.4]
  assign storesToCheck_1_3 = _T_1346 ? _T_3473 : _T_3480; // @[LoadQueue.scala 131:10:@3513.4]
  assign _T_3486 = 3'h4 <= offsetQ_1; // @[LoadQueue.scala 131:81:@3516.4]
  assign _T_3487 = _T_2855 & _T_3486; // @[LoadQueue.scala 131:72:@3517.4]
  assign _T_3489 = offsetQ_1 < 3'h4; // @[LoadQueue.scala 132:33:@3518.4]
  assign _T_3492 = _T_3489 & _T_2864; // @[LoadQueue.scala 132:41:@3520.4]
  assign _T_3494 = _T_3492 == 1'h0; // @[LoadQueue.scala 132:9:@3521.4]
  assign storesToCheck_1_4 = _T_1346 ? _T_3487 : _T_3494; // @[LoadQueue.scala 131:10:@3522.4]
  assign _T_3500 = 3'h5 <= offsetQ_1; // @[LoadQueue.scala 131:81:@3525.4]
  assign _T_3501 = _T_2872 & _T_3500; // @[LoadQueue.scala 131:72:@3526.4]
  assign _T_3503 = offsetQ_1 < 3'h5; // @[LoadQueue.scala 132:33:@3527.4]
  assign _T_3506 = _T_3503 & _T_2881; // @[LoadQueue.scala 132:41:@3529.4]
  assign _T_3508 = _T_3506 == 1'h0; // @[LoadQueue.scala 132:9:@3530.4]
  assign storesToCheck_1_5 = _T_1346 ? _T_3501 : _T_3508; // @[LoadQueue.scala 131:10:@3531.4]
  assign _T_3514 = 3'h6 <= offsetQ_1; // @[LoadQueue.scala 131:81:@3534.4]
  assign _T_3515 = _T_2889 & _T_3514; // @[LoadQueue.scala 131:72:@3535.4]
  assign _T_3517 = offsetQ_1 < 3'h6; // @[LoadQueue.scala 132:33:@3536.4]
  assign _T_3520 = _T_3517 & _T_2898; // @[LoadQueue.scala 132:41:@3538.4]
  assign _T_3522 = _T_3520 == 1'h0; // @[LoadQueue.scala 132:9:@3539.4]
  assign storesToCheck_1_6 = _T_1346 ? _T_3515 : _T_3522; // @[LoadQueue.scala 131:10:@3540.4]
  assign _T_3528 = 3'h7 <= offsetQ_1; // @[LoadQueue.scala 131:81:@3543.4]
  assign storesToCheck_1_7 = _T_1346 ? _T_3528 : 1'h1; // @[LoadQueue.scala 131:10:@3549.4]
  assign storesToCheck_2_0 = _T_1376 ? _T_2787 : 1'h1; // @[LoadQueue.scala 131:10:@3575.4]
  assign _T_3570 = 3'h1 <= offsetQ_2; // @[LoadQueue.scala 131:81:@3578.4]
  assign _T_3571 = _T_2804 & _T_3570; // @[LoadQueue.scala 131:72:@3579.4]
  assign _T_3573 = offsetQ_2 < 3'h1; // @[LoadQueue.scala 132:33:@3580.4]
  assign _T_3576 = _T_3573 & _T_2813; // @[LoadQueue.scala 132:41:@3582.4]
  assign _T_3578 = _T_3576 == 1'h0; // @[LoadQueue.scala 132:9:@3583.4]
  assign storesToCheck_2_1 = _T_1376 ? _T_3571 : _T_3578; // @[LoadQueue.scala 131:10:@3584.4]
  assign _T_3584 = 3'h2 <= offsetQ_2; // @[LoadQueue.scala 131:81:@3587.4]
  assign _T_3585 = _T_2821 & _T_3584; // @[LoadQueue.scala 131:72:@3588.4]
  assign _T_3587 = offsetQ_2 < 3'h2; // @[LoadQueue.scala 132:33:@3589.4]
  assign _T_3590 = _T_3587 & _T_2830; // @[LoadQueue.scala 132:41:@3591.4]
  assign _T_3592 = _T_3590 == 1'h0; // @[LoadQueue.scala 132:9:@3592.4]
  assign storesToCheck_2_2 = _T_1376 ? _T_3585 : _T_3592; // @[LoadQueue.scala 131:10:@3593.4]
  assign _T_3598 = 3'h3 <= offsetQ_2; // @[LoadQueue.scala 131:81:@3596.4]
  assign _T_3599 = _T_2838 & _T_3598; // @[LoadQueue.scala 131:72:@3597.4]
  assign _T_3601 = offsetQ_2 < 3'h3; // @[LoadQueue.scala 132:33:@3598.4]
  assign _T_3604 = _T_3601 & _T_2847; // @[LoadQueue.scala 132:41:@3600.4]
  assign _T_3606 = _T_3604 == 1'h0; // @[LoadQueue.scala 132:9:@3601.4]
  assign storesToCheck_2_3 = _T_1376 ? _T_3599 : _T_3606; // @[LoadQueue.scala 131:10:@3602.4]
  assign _T_3612 = 3'h4 <= offsetQ_2; // @[LoadQueue.scala 131:81:@3605.4]
  assign _T_3613 = _T_2855 & _T_3612; // @[LoadQueue.scala 131:72:@3606.4]
  assign _T_3615 = offsetQ_2 < 3'h4; // @[LoadQueue.scala 132:33:@3607.4]
  assign _T_3618 = _T_3615 & _T_2864; // @[LoadQueue.scala 132:41:@3609.4]
  assign _T_3620 = _T_3618 == 1'h0; // @[LoadQueue.scala 132:9:@3610.4]
  assign storesToCheck_2_4 = _T_1376 ? _T_3613 : _T_3620; // @[LoadQueue.scala 131:10:@3611.4]
  assign _T_3626 = 3'h5 <= offsetQ_2; // @[LoadQueue.scala 131:81:@3614.4]
  assign _T_3627 = _T_2872 & _T_3626; // @[LoadQueue.scala 131:72:@3615.4]
  assign _T_3629 = offsetQ_2 < 3'h5; // @[LoadQueue.scala 132:33:@3616.4]
  assign _T_3632 = _T_3629 & _T_2881; // @[LoadQueue.scala 132:41:@3618.4]
  assign _T_3634 = _T_3632 == 1'h0; // @[LoadQueue.scala 132:9:@3619.4]
  assign storesToCheck_2_5 = _T_1376 ? _T_3627 : _T_3634; // @[LoadQueue.scala 131:10:@3620.4]
  assign _T_3640 = 3'h6 <= offsetQ_2; // @[LoadQueue.scala 131:81:@3623.4]
  assign _T_3641 = _T_2889 & _T_3640; // @[LoadQueue.scala 131:72:@3624.4]
  assign _T_3643 = offsetQ_2 < 3'h6; // @[LoadQueue.scala 132:33:@3625.4]
  assign _T_3646 = _T_3643 & _T_2898; // @[LoadQueue.scala 132:41:@3627.4]
  assign _T_3648 = _T_3646 == 1'h0; // @[LoadQueue.scala 132:9:@3628.4]
  assign storesToCheck_2_6 = _T_1376 ? _T_3641 : _T_3648; // @[LoadQueue.scala 131:10:@3629.4]
  assign _T_3654 = 3'h7 <= offsetQ_2; // @[LoadQueue.scala 131:81:@3632.4]
  assign storesToCheck_2_7 = _T_1376 ? _T_3654 : 1'h1; // @[LoadQueue.scala 131:10:@3638.4]
  assign storesToCheck_3_0 = _T_1406 ? _T_2787 : 1'h1; // @[LoadQueue.scala 131:10:@3664.4]
  assign _T_3696 = 3'h1 <= offsetQ_3; // @[LoadQueue.scala 131:81:@3667.4]
  assign _T_3697 = _T_2804 & _T_3696; // @[LoadQueue.scala 131:72:@3668.4]
  assign _T_3699 = offsetQ_3 < 3'h1; // @[LoadQueue.scala 132:33:@3669.4]
  assign _T_3702 = _T_3699 & _T_2813; // @[LoadQueue.scala 132:41:@3671.4]
  assign _T_3704 = _T_3702 == 1'h0; // @[LoadQueue.scala 132:9:@3672.4]
  assign storesToCheck_3_1 = _T_1406 ? _T_3697 : _T_3704; // @[LoadQueue.scala 131:10:@3673.4]
  assign _T_3710 = 3'h2 <= offsetQ_3; // @[LoadQueue.scala 131:81:@3676.4]
  assign _T_3711 = _T_2821 & _T_3710; // @[LoadQueue.scala 131:72:@3677.4]
  assign _T_3713 = offsetQ_3 < 3'h2; // @[LoadQueue.scala 132:33:@3678.4]
  assign _T_3716 = _T_3713 & _T_2830; // @[LoadQueue.scala 132:41:@3680.4]
  assign _T_3718 = _T_3716 == 1'h0; // @[LoadQueue.scala 132:9:@3681.4]
  assign storesToCheck_3_2 = _T_1406 ? _T_3711 : _T_3718; // @[LoadQueue.scala 131:10:@3682.4]
  assign _T_3724 = 3'h3 <= offsetQ_3; // @[LoadQueue.scala 131:81:@3685.4]
  assign _T_3725 = _T_2838 & _T_3724; // @[LoadQueue.scala 131:72:@3686.4]
  assign _T_3727 = offsetQ_3 < 3'h3; // @[LoadQueue.scala 132:33:@3687.4]
  assign _T_3730 = _T_3727 & _T_2847; // @[LoadQueue.scala 132:41:@3689.4]
  assign _T_3732 = _T_3730 == 1'h0; // @[LoadQueue.scala 132:9:@3690.4]
  assign storesToCheck_3_3 = _T_1406 ? _T_3725 : _T_3732; // @[LoadQueue.scala 131:10:@3691.4]
  assign _T_3738 = 3'h4 <= offsetQ_3; // @[LoadQueue.scala 131:81:@3694.4]
  assign _T_3739 = _T_2855 & _T_3738; // @[LoadQueue.scala 131:72:@3695.4]
  assign _T_3741 = offsetQ_3 < 3'h4; // @[LoadQueue.scala 132:33:@3696.4]
  assign _T_3744 = _T_3741 & _T_2864; // @[LoadQueue.scala 132:41:@3698.4]
  assign _T_3746 = _T_3744 == 1'h0; // @[LoadQueue.scala 132:9:@3699.4]
  assign storesToCheck_3_4 = _T_1406 ? _T_3739 : _T_3746; // @[LoadQueue.scala 131:10:@3700.4]
  assign _T_3752 = 3'h5 <= offsetQ_3; // @[LoadQueue.scala 131:81:@3703.4]
  assign _T_3753 = _T_2872 & _T_3752; // @[LoadQueue.scala 131:72:@3704.4]
  assign _T_3755 = offsetQ_3 < 3'h5; // @[LoadQueue.scala 132:33:@3705.4]
  assign _T_3758 = _T_3755 & _T_2881; // @[LoadQueue.scala 132:41:@3707.4]
  assign _T_3760 = _T_3758 == 1'h0; // @[LoadQueue.scala 132:9:@3708.4]
  assign storesToCheck_3_5 = _T_1406 ? _T_3753 : _T_3760; // @[LoadQueue.scala 131:10:@3709.4]
  assign _T_3766 = 3'h6 <= offsetQ_3; // @[LoadQueue.scala 131:81:@3712.4]
  assign _T_3767 = _T_2889 & _T_3766; // @[LoadQueue.scala 131:72:@3713.4]
  assign _T_3769 = offsetQ_3 < 3'h6; // @[LoadQueue.scala 132:33:@3714.4]
  assign _T_3772 = _T_3769 & _T_2898; // @[LoadQueue.scala 132:41:@3716.4]
  assign _T_3774 = _T_3772 == 1'h0; // @[LoadQueue.scala 132:9:@3717.4]
  assign storesToCheck_3_6 = _T_1406 ? _T_3767 : _T_3774; // @[LoadQueue.scala 131:10:@3718.4]
  assign _T_3780 = 3'h7 <= offsetQ_3; // @[LoadQueue.scala 131:81:@3721.4]
  assign storesToCheck_3_7 = _T_1406 ? _T_3780 : 1'h1; // @[LoadQueue.scala 131:10:@3727.4]
  assign storesToCheck_4_0 = _T_1436 ? _T_2787 : 1'h1; // @[LoadQueue.scala 131:10:@3753.4]
  assign _T_3822 = 3'h1 <= offsetQ_4; // @[LoadQueue.scala 131:81:@3756.4]
  assign _T_3823 = _T_2804 & _T_3822; // @[LoadQueue.scala 131:72:@3757.4]
  assign _T_3825 = offsetQ_4 < 3'h1; // @[LoadQueue.scala 132:33:@3758.4]
  assign _T_3828 = _T_3825 & _T_2813; // @[LoadQueue.scala 132:41:@3760.4]
  assign _T_3830 = _T_3828 == 1'h0; // @[LoadQueue.scala 132:9:@3761.4]
  assign storesToCheck_4_1 = _T_1436 ? _T_3823 : _T_3830; // @[LoadQueue.scala 131:10:@3762.4]
  assign _T_3836 = 3'h2 <= offsetQ_4; // @[LoadQueue.scala 131:81:@3765.4]
  assign _T_3837 = _T_2821 & _T_3836; // @[LoadQueue.scala 131:72:@3766.4]
  assign _T_3839 = offsetQ_4 < 3'h2; // @[LoadQueue.scala 132:33:@3767.4]
  assign _T_3842 = _T_3839 & _T_2830; // @[LoadQueue.scala 132:41:@3769.4]
  assign _T_3844 = _T_3842 == 1'h0; // @[LoadQueue.scala 132:9:@3770.4]
  assign storesToCheck_4_2 = _T_1436 ? _T_3837 : _T_3844; // @[LoadQueue.scala 131:10:@3771.4]
  assign _T_3850 = 3'h3 <= offsetQ_4; // @[LoadQueue.scala 131:81:@3774.4]
  assign _T_3851 = _T_2838 & _T_3850; // @[LoadQueue.scala 131:72:@3775.4]
  assign _T_3853 = offsetQ_4 < 3'h3; // @[LoadQueue.scala 132:33:@3776.4]
  assign _T_3856 = _T_3853 & _T_2847; // @[LoadQueue.scala 132:41:@3778.4]
  assign _T_3858 = _T_3856 == 1'h0; // @[LoadQueue.scala 132:9:@3779.4]
  assign storesToCheck_4_3 = _T_1436 ? _T_3851 : _T_3858; // @[LoadQueue.scala 131:10:@3780.4]
  assign _T_3864 = 3'h4 <= offsetQ_4; // @[LoadQueue.scala 131:81:@3783.4]
  assign _T_3865 = _T_2855 & _T_3864; // @[LoadQueue.scala 131:72:@3784.4]
  assign _T_3867 = offsetQ_4 < 3'h4; // @[LoadQueue.scala 132:33:@3785.4]
  assign _T_3870 = _T_3867 & _T_2864; // @[LoadQueue.scala 132:41:@3787.4]
  assign _T_3872 = _T_3870 == 1'h0; // @[LoadQueue.scala 132:9:@3788.4]
  assign storesToCheck_4_4 = _T_1436 ? _T_3865 : _T_3872; // @[LoadQueue.scala 131:10:@3789.4]
  assign _T_3878 = 3'h5 <= offsetQ_4; // @[LoadQueue.scala 131:81:@3792.4]
  assign _T_3879 = _T_2872 & _T_3878; // @[LoadQueue.scala 131:72:@3793.4]
  assign _T_3881 = offsetQ_4 < 3'h5; // @[LoadQueue.scala 132:33:@3794.4]
  assign _T_3884 = _T_3881 & _T_2881; // @[LoadQueue.scala 132:41:@3796.4]
  assign _T_3886 = _T_3884 == 1'h0; // @[LoadQueue.scala 132:9:@3797.4]
  assign storesToCheck_4_5 = _T_1436 ? _T_3879 : _T_3886; // @[LoadQueue.scala 131:10:@3798.4]
  assign _T_3892 = 3'h6 <= offsetQ_4; // @[LoadQueue.scala 131:81:@3801.4]
  assign _T_3893 = _T_2889 & _T_3892; // @[LoadQueue.scala 131:72:@3802.4]
  assign _T_3895 = offsetQ_4 < 3'h6; // @[LoadQueue.scala 132:33:@3803.4]
  assign _T_3898 = _T_3895 & _T_2898; // @[LoadQueue.scala 132:41:@3805.4]
  assign _T_3900 = _T_3898 == 1'h0; // @[LoadQueue.scala 132:9:@3806.4]
  assign storesToCheck_4_6 = _T_1436 ? _T_3893 : _T_3900; // @[LoadQueue.scala 131:10:@3807.4]
  assign _T_3906 = 3'h7 <= offsetQ_4; // @[LoadQueue.scala 131:81:@3810.4]
  assign storesToCheck_4_7 = _T_1436 ? _T_3906 : 1'h1; // @[LoadQueue.scala 131:10:@3816.4]
  assign storesToCheck_5_0 = _T_1466 ? _T_2787 : 1'h1; // @[LoadQueue.scala 131:10:@3842.4]
  assign _T_3948 = 3'h1 <= offsetQ_5; // @[LoadQueue.scala 131:81:@3845.4]
  assign _T_3949 = _T_2804 & _T_3948; // @[LoadQueue.scala 131:72:@3846.4]
  assign _T_3951 = offsetQ_5 < 3'h1; // @[LoadQueue.scala 132:33:@3847.4]
  assign _T_3954 = _T_3951 & _T_2813; // @[LoadQueue.scala 132:41:@3849.4]
  assign _T_3956 = _T_3954 == 1'h0; // @[LoadQueue.scala 132:9:@3850.4]
  assign storesToCheck_5_1 = _T_1466 ? _T_3949 : _T_3956; // @[LoadQueue.scala 131:10:@3851.4]
  assign _T_3962 = 3'h2 <= offsetQ_5; // @[LoadQueue.scala 131:81:@3854.4]
  assign _T_3963 = _T_2821 & _T_3962; // @[LoadQueue.scala 131:72:@3855.4]
  assign _T_3965 = offsetQ_5 < 3'h2; // @[LoadQueue.scala 132:33:@3856.4]
  assign _T_3968 = _T_3965 & _T_2830; // @[LoadQueue.scala 132:41:@3858.4]
  assign _T_3970 = _T_3968 == 1'h0; // @[LoadQueue.scala 132:9:@3859.4]
  assign storesToCheck_5_2 = _T_1466 ? _T_3963 : _T_3970; // @[LoadQueue.scala 131:10:@3860.4]
  assign _T_3976 = 3'h3 <= offsetQ_5; // @[LoadQueue.scala 131:81:@3863.4]
  assign _T_3977 = _T_2838 & _T_3976; // @[LoadQueue.scala 131:72:@3864.4]
  assign _T_3979 = offsetQ_5 < 3'h3; // @[LoadQueue.scala 132:33:@3865.4]
  assign _T_3982 = _T_3979 & _T_2847; // @[LoadQueue.scala 132:41:@3867.4]
  assign _T_3984 = _T_3982 == 1'h0; // @[LoadQueue.scala 132:9:@3868.4]
  assign storesToCheck_5_3 = _T_1466 ? _T_3977 : _T_3984; // @[LoadQueue.scala 131:10:@3869.4]
  assign _T_3990 = 3'h4 <= offsetQ_5; // @[LoadQueue.scala 131:81:@3872.4]
  assign _T_3991 = _T_2855 & _T_3990; // @[LoadQueue.scala 131:72:@3873.4]
  assign _T_3993 = offsetQ_5 < 3'h4; // @[LoadQueue.scala 132:33:@3874.4]
  assign _T_3996 = _T_3993 & _T_2864; // @[LoadQueue.scala 132:41:@3876.4]
  assign _T_3998 = _T_3996 == 1'h0; // @[LoadQueue.scala 132:9:@3877.4]
  assign storesToCheck_5_4 = _T_1466 ? _T_3991 : _T_3998; // @[LoadQueue.scala 131:10:@3878.4]
  assign _T_4004 = 3'h5 <= offsetQ_5; // @[LoadQueue.scala 131:81:@3881.4]
  assign _T_4005 = _T_2872 & _T_4004; // @[LoadQueue.scala 131:72:@3882.4]
  assign _T_4007 = offsetQ_5 < 3'h5; // @[LoadQueue.scala 132:33:@3883.4]
  assign _T_4010 = _T_4007 & _T_2881; // @[LoadQueue.scala 132:41:@3885.4]
  assign _T_4012 = _T_4010 == 1'h0; // @[LoadQueue.scala 132:9:@3886.4]
  assign storesToCheck_5_5 = _T_1466 ? _T_4005 : _T_4012; // @[LoadQueue.scala 131:10:@3887.4]
  assign _T_4018 = 3'h6 <= offsetQ_5; // @[LoadQueue.scala 131:81:@3890.4]
  assign _T_4019 = _T_2889 & _T_4018; // @[LoadQueue.scala 131:72:@3891.4]
  assign _T_4021 = offsetQ_5 < 3'h6; // @[LoadQueue.scala 132:33:@3892.4]
  assign _T_4024 = _T_4021 & _T_2898; // @[LoadQueue.scala 132:41:@3894.4]
  assign _T_4026 = _T_4024 == 1'h0; // @[LoadQueue.scala 132:9:@3895.4]
  assign storesToCheck_5_6 = _T_1466 ? _T_4019 : _T_4026; // @[LoadQueue.scala 131:10:@3896.4]
  assign _T_4032 = 3'h7 <= offsetQ_5; // @[LoadQueue.scala 131:81:@3899.4]
  assign storesToCheck_5_7 = _T_1466 ? _T_4032 : 1'h1; // @[LoadQueue.scala 131:10:@3905.4]
  assign storesToCheck_6_0 = _T_1496 ? _T_2787 : 1'h1; // @[LoadQueue.scala 131:10:@3931.4]
  assign _T_4074 = 3'h1 <= offsetQ_6; // @[LoadQueue.scala 131:81:@3934.4]
  assign _T_4075 = _T_2804 & _T_4074; // @[LoadQueue.scala 131:72:@3935.4]
  assign _T_4077 = offsetQ_6 < 3'h1; // @[LoadQueue.scala 132:33:@3936.4]
  assign _T_4080 = _T_4077 & _T_2813; // @[LoadQueue.scala 132:41:@3938.4]
  assign _T_4082 = _T_4080 == 1'h0; // @[LoadQueue.scala 132:9:@3939.4]
  assign storesToCheck_6_1 = _T_1496 ? _T_4075 : _T_4082; // @[LoadQueue.scala 131:10:@3940.4]
  assign _T_4088 = 3'h2 <= offsetQ_6; // @[LoadQueue.scala 131:81:@3943.4]
  assign _T_4089 = _T_2821 & _T_4088; // @[LoadQueue.scala 131:72:@3944.4]
  assign _T_4091 = offsetQ_6 < 3'h2; // @[LoadQueue.scala 132:33:@3945.4]
  assign _T_4094 = _T_4091 & _T_2830; // @[LoadQueue.scala 132:41:@3947.4]
  assign _T_4096 = _T_4094 == 1'h0; // @[LoadQueue.scala 132:9:@3948.4]
  assign storesToCheck_6_2 = _T_1496 ? _T_4089 : _T_4096; // @[LoadQueue.scala 131:10:@3949.4]
  assign _T_4102 = 3'h3 <= offsetQ_6; // @[LoadQueue.scala 131:81:@3952.4]
  assign _T_4103 = _T_2838 & _T_4102; // @[LoadQueue.scala 131:72:@3953.4]
  assign _T_4105 = offsetQ_6 < 3'h3; // @[LoadQueue.scala 132:33:@3954.4]
  assign _T_4108 = _T_4105 & _T_2847; // @[LoadQueue.scala 132:41:@3956.4]
  assign _T_4110 = _T_4108 == 1'h0; // @[LoadQueue.scala 132:9:@3957.4]
  assign storesToCheck_6_3 = _T_1496 ? _T_4103 : _T_4110; // @[LoadQueue.scala 131:10:@3958.4]
  assign _T_4116 = 3'h4 <= offsetQ_6; // @[LoadQueue.scala 131:81:@3961.4]
  assign _T_4117 = _T_2855 & _T_4116; // @[LoadQueue.scala 131:72:@3962.4]
  assign _T_4119 = offsetQ_6 < 3'h4; // @[LoadQueue.scala 132:33:@3963.4]
  assign _T_4122 = _T_4119 & _T_2864; // @[LoadQueue.scala 132:41:@3965.4]
  assign _T_4124 = _T_4122 == 1'h0; // @[LoadQueue.scala 132:9:@3966.4]
  assign storesToCheck_6_4 = _T_1496 ? _T_4117 : _T_4124; // @[LoadQueue.scala 131:10:@3967.4]
  assign _T_4130 = 3'h5 <= offsetQ_6; // @[LoadQueue.scala 131:81:@3970.4]
  assign _T_4131 = _T_2872 & _T_4130; // @[LoadQueue.scala 131:72:@3971.4]
  assign _T_4133 = offsetQ_6 < 3'h5; // @[LoadQueue.scala 132:33:@3972.4]
  assign _T_4136 = _T_4133 & _T_2881; // @[LoadQueue.scala 132:41:@3974.4]
  assign _T_4138 = _T_4136 == 1'h0; // @[LoadQueue.scala 132:9:@3975.4]
  assign storesToCheck_6_5 = _T_1496 ? _T_4131 : _T_4138; // @[LoadQueue.scala 131:10:@3976.4]
  assign _T_4144 = 3'h6 <= offsetQ_6; // @[LoadQueue.scala 131:81:@3979.4]
  assign _T_4145 = _T_2889 & _T_4144; // @[LoadQueue.scala 131:72:@3980.4]
  assign _T_4147 = offsetQ_6 < 3'h6; // @[LoadQueue.scala 132:33:@3981.4]
  assign _T_4150 = _T_4147 & _T_2898; // @[LoadQueue.scala 132:41:@3983.4]
  assign _T_4152 = _T_4150 == 1'h0; // @[LoadQueue.scala 132:9:@3984.4]
  assign storesToCheck_6_6 = _T_1496 ? _T_4145 : _T_4152; // @[LoadQueue.scala 131:10:@3985.4]
  assign _T_4158 = 3'h7 <= offsetQ_6; // @[LoadQueue.scala 131:81:@3988.4]
  assign storesToCheck_6_7 = _T_1496 ? _T_4158 : 1'h1; // @[LoadQueue.scala 131:10:@3994.4]
  assign storesToCheck_7_0 = _T_1526 ? _T_2787 : 1'h1; // @[LoadQueue.scala 131:10:@4020.4]
  assign _T_4200 = 3'h1 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4023.4]
  assign _T_4201 = _T_2804 & _T_4200; // @[LoadQueue.scala 131:72:@4024.4]
  assign _T_4203 = offsetQ_7 < 3'h1; // @[LoadQueue.scala 132:33:@4025.4]
  assign _T_4206 = _T_4203 & _T_2813; // @[LoadQueue.scala 132:41:@4027.4]
  assign _T_4208 = _T_4206 == 1'h0; // @[LoadQueue.scala 132:9:@4028.4]
  assign storesToCheck_7_1 = _T_1526 ? _T_4201 : _T_4208; // @[LoadQueue.scala 131:10:@4029.4]
  assign _T_4214 = 3'h2 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4032.4]
  assign _T_4215 = _T_2821 & _T_4214; // @[LoadQueue.scala 131:72:@4033.4]
  assign _T_4217 = offsetQ_7 < 3'h2; // @[LoadQueue.scala 132:33:@4034.4]
  assign _T_4220 = _T_4217 & _T_2830; // @[LoadQueue.scala 132:41:@4036.4]
  assign _T_4222 = _T_4220 == 1'h0; // @[LoadQueue.scala 132:9:@4037.4]
  assign storesToCheck_7_2 = _T_1526 ? _T_4215 : _T_4222; // @[LoadQueue.scala 131:10:@4038.4]
  assign _T_4228 = 3'h3 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4041.4]
  assign _T_4229 = _T_2838 & _T_4228; // @[LoadQueue.scala 131:72:@4042.4]
  assign _T_4231 = offsetQ_7 < 3'h3; // @[LoadQueue.scala 132:33:@4043.4]
  assign _T_4234 = _T_4231 & _T_2847; // @[LoadQueue.scala 132:41:@4045.4]
  assign _T_4236 = _T_4234 == 1'h0; // @[LoadQueue.scala 132:9:@4046.4]
  assign storesToCheck_7_3 = _T_1526 ? _T_4229 : _T_4236; // @[LoadQueue.scala 131:10:@4047.4]
  assign _T_4242 = 3'h4 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4050.4]
  assign _T_4243 = _T_2855 & _T_4242; // @[LoadQueue.scala 131:72:@4051.4]
  assign _T_4245 = offsetQ_7 < 3'h4; // @[LoadQueue.scala 132:33:@4052.4]
  assign _T_4248 = _T_4245 & _T_2864; // @[LoadQueue.scala 132:41:@4054.4]
  assign _T_4250 = _T_4248 == 1'h0; // @[LoadQueue.scala 132:9:@4055.4]
  assign storesToCheck_7_4 = _T_1526 ? _T_4243 : _T_4250; // @[LoadQueue.scala 131:10:@4056.4]
  assign _T_4256 = 3'h5 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4059.4]
  assign _T_4257 = _T_2872 & _T_4256; // @[LoadQueue.scala 131:72:@4060.4]
  assign _T_4259 = offsetQ_7 < 3'h5; // @[LoadQueue.scala 132:33:@4061.4]
  assign _T_4262 = _T_4259 & _T_2881; // @[LoadQueue.scala 132:41:@4063.4]
  assign _T_4264 = _T_4262 == 1'h0; // @[LoadQueue.scala 132:9:@4064.4]
  assign storesToCheck_7_5 = _T_1526 ? _T_4257 : _T_4264; // @[LoadQueue.scala 131:10:@4065.4]
  assign _T_4270 = 3'h6 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4068.4]
  assign _T_4271 = _T_2889 & _T_4270; // @[LoadQueue.scala 131:72:@4069.4]
  assign _T_4273 = offsetQ_7 < 3'h6; // @[LoadQueue.scala 132:33:@4070.4]
  assign _T_4276 = _T_4273 & _T_2898; // @[LoadQueue.scala 132:41:@4072.4]
  assign _T_4278 = _T_4276 == 1'h0; // @[LoadQueue.scala 132:9:@4073.4]
  assign storesToCheck_7_6 = _T_1526 ? _T_4271 : _T_4278; // @[LoadQueue.scala 131:10:@4074.4]
  assign _T_4284 = 3'h7 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4077.4]
  assign storesToCheck_7_7 = _T_1526 ? _T_4284 : 1'h1; // @[LoadQueue.scala 131:10:@4083.4]
  assign _T_4674 = storesToCheck_0_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4102.4]
  assign entriesToCheck_0_0 = _T_4674 & checkBits_0; // @[LoadQueue.scala 141:26:@4103.4]
  assign _T_4676 = storesToCheck_0_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4104.4]
  assign entriesToCheck_0_1 = _T_4676 & checkBits_0; // @[LoadQueue.scala 141:26:@4105.4]
  assign _T_4678 = storesToCheck_0_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4106.4]
  assign entriesToCheck_0_2 = _T_4678 & checkBits_0; // @[LoadQueue.scala 141:26:@4107.4]
  assign _T_4680 = storesToCheck_0_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4108.4]
  assign entriesToCheck_0_3 = _T_4680 & checkBits_0; // @[LoadQueue.scala 141:26:@4109.4]
  assign _T_4682 = storesToCheck_0_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4110.4]
  assign entriesToCheck_0_4 = _T_4682 & checkBits_0; // @[LoadQueue.scala 141:26:@4111.4]
  assign _T_4684 = storesToCheck_0_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4112.4]
  assign entriesToCheck_0_5 = _T_4684 & checkBits_0; // @[LoadQueue.scala 141:26:@4113.4]
  assign _T_4686 = storesToCheck_0_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4114.4]
  assign entriesToCheck_0_6 = _T_4686 & checkBits_0; // @[LoadQueue.scala 141:26:@4115.4]
  assign _T_4688 = storesToCheck_0_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4116.4]
  assign entriesToCheck_0_7 = _T_4688 & checkBits_0; // @[LoadQueue.scala 141:26:@4117.4]
  assign _T_4690 = storesToCheck_1_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4126.4]
  assign entriesToCheck_1_0 = _T_4690 & checkBits_1; // @[LoadQueue.scala 141:26:@4127.4]
  assign _T_4692 = storesToCheck_1_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4128.4]
  assign entriesToCheck_1_1 = _T_4692 & checkBits_1; // @[LoadQueue.scala 141:26:@4129.4]
  assign _T_4694 = storesToCheck_1_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4130.4]
  assign entriesToCheck_1_2 = _T_4694 & checkBits_1; // @[LoadQueue.scala 141:26:@4131.4]
  assign _T_4696 = storesToCheck_1_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4132.4]
  assign entriesToCheck_1_3 = _T_4696 & checkBits_1; // @[LoadQueue.scala 141:26:@4133.4]
  assign _T_4698 = storesToCheck_1_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4134.4]
  assign entriesToCheck_1_4 = _T_4698 & checkBits_1; // @[LoadQueue.scala 141:26:@4135.4]
  assign _T_4700 = storesToCheck_1_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4136.4]
  assign entriesToCheck_1_5 = _T_4700 & checkBits_1; // @[LoadQueue.scala 141:26:@4137.4]
  assign _T_4702 = storesToCheck_1_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4138.4]
  assign entriesToCheck_1_6 = _T_4702 & checkBits_1; // @[LoadQueue.scala 141:26:@4139.4]
  assign _T_4704 = storesToCheck_1_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4140.4]
  assign entriesToCheck_1_7 = _T_4704 & checkBits_1; // @[LoadQueue.scala 141:26:@4141.4]
  assign _T_4706 = storesToCheck_2_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4150.4]
  assign entriesToCheck_2_0 = _T_4706 & checkBits_2; // @[LoadQueue.scala 141:26:@4151.4]
  assign _T_4708 = storesToCheck_2_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4152.4]
  assign entriesToCheck_2_1 = _T_4708 & checkBits_2; // @[LoadQueue.scala 141:26:@4153.4]
  assign _T_4710 = storesToCheck_2_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4154.4]
  assign entriesToCheck_2_2 = _T_4710 & checkBits_2; // @[LoadQueue.scala 141:26:@4155.4]
  assign _T_4712 = storesToCheck_2_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4156.4]
  assign entriesToCheck_2_3 = _T_4712 & checkBits_2; // @[LoadQueue.scala 141:26:@4157.4]
  assign _T_4714 = storesToCheck_2_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4158.4]
  assign entriesToCheck_2_4 = _T_4714 & checkBits_2; // @[LoadQueue.scala 141:26:@4159.4]
  assign _T_4716 = storesToCheck_2_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4160.4]
  assign entriesToCheck_2_5 = _T_4716 & checkBits_2; // @[LoadQueue.scala 141:26:@4161.4]
  assign _T_4718 = storesToCheck_2_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4162.4]
  assign entriesToCheck_2_6 = _T_4718 & checkBits_2; // @[LoadQueue.scala 141:26:@4163.4]
  assign _T_4720 = storesToCheck_2_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4164.4]
  assign entriesToCheck_2_7 = _T_4720 & checkBits_2; // @[LoadQueue.scala 141:26:@4165.4]
  assign _T_4722 = storesToCheck_3_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4174.4]
  assign entriesToCheck_3_0 = _T_4722 & checkBits_3; // @[LoadQueue.scala 141:26:@4175.4]
  assign _T_4724 = storesToCheck_3_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4176.4]
  assign entriesToCheck_3_1 = _T_4724 & checkBits_3; // @[LoadQueue.scala 141:26:@4177.4]
  assign _T_4726 = storesToCheck_3_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4178.4]
  assign entriesToCheck_3_2 = _T_4726 & checkBits_3; // @[LoadQueue.scala 141:26:@4179.4]
  assign _T_4728 = storesToCheck_3_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4180.4]
  assign entriesToCheck_3_3 = _T_4728 & checkBits_3; // @[LoadQueue.scala 141:26:@4181.4]
  assign _T_4730 = storesToCheck_3_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4182.4]
  assign entriesToCheck_3_4 = _T_4730 & checkBits_3; // @[LoadQueue.scala 141:26:@4183.4]
  assign _T_4732 = storesToCheck_3_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4184.4]
  assign entriesToCheck_3_5 = _T_4732 & checkBits_3; // @[LoadQueue.scala 141:26:@4185.4]
  assign _T_4734 = storesToCheck_3_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4186.4]
  assign entriesToCheck_3_6 = _T_4734 & checkBits_3; // @[LoadQueue.scala 141:26:@4187.4]
  assign _T_4736 = storesToCheck_3_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4188.4]
  assign entriesToCheck_3_7 = _T_4736 & checkBits_3; // @[LoadQueue.scala 141:26:@4189.4]
  assign _T_4738 = storesToCheck_4_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4198.4]
  assign entriesToCheck_4_0 = _T_4738 & checkBits_4; // @[LoadQueue.scala 141:26:@4199.4]
  assign _T_4740 = storesToCheck_4_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4200.4]
  assign entriesToCheck_4_1 = _T_4740 & checkBits_4; // @[LoadQueue.scala 141:26:@4201.4]
  assign _T_4742 = storesToCheck_4_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4202.4]
  assign entriesToCheck_4_2 = _T_4742 & checkBits_4; // @[LoadQueue.scala 141:26:@4203.4]
  assign _T_4744 = storesToCheck_4_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4204.4]
  assign entriesToCheck_4_3 = _T_4744 & checkBits_4; // @[LoadQueue.scala 141:26:@4205.4]
  assign _T_4746 = storesToCheck_4_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4206.4]
  assign entriesToCheck_4_4 = _T_4746 & checkBits_4; // @[LoadQueue.scala 141:26:@4207.4]
  assign _T_4748 = storesToCheck_4_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4208.4]
  assign entriesToCheck_4_5 = _T_4748 & checkBits_4; // @[LoadQueue.scala 141:26:@4209.4]
  assign _T_4750 = storesToCheck_4_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4210.4]
  assign entriesToCheck_4_6 = _T_4750 & checkBits_4; // @[LoadQueue.scala 141:26:@4211.4]
  assign _T_4752 = storesToCheck_4_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4212.4]
  assign entriesToCheck_4_7 = _T_4752 & checkBits_4; // @[LoadQueue.scala 141:26:@4213.4]
  assign _T_4754 = storesToCheck_5_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4222.4]
  assign entriesToCheck_5_0 = _T_4754 & checkBits_5; // @[LoadQueue.scala 141:26:@4223.4]
  assign _T_4756 = storesToCheck_5_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4224.4]
  assign entriesToCheck_5_1 = _T_4756 & checkBits_5; // @[LoadQueue.scala 141:26:@4225.4]
  assign _T_4758 = storesToCheck_5_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4226.4]
  assign entriesToCheck_5_2 = _T_4758 & checkBits_5; // @[LoadQueue.scala 141:26:@4227.4]
  assign _T_4760 = storesToCheck_5_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4228.4]
  assign entriesToCheck_5_3 = _T_4760 & checkBits_5; // @[LoadQueue.scala 141:26:@4229.4]
  assign _T_4762 = storesToCheck_5_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4230.4]
  assign entriesToCheck_5_4 = _T_4762 & checkBits_5; // @[LoadQueue.scala 141:26:@4231.4]
  assign _T_4764 = storesToCheck_5_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4232.4]
  assign entriesToCheck_5_5 = _T_4764 & checkBits_5; // @[LoadQueue.scala 141:26:@4233.4]
  assign _T_4766 = storesToCheck_5_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4234.4]
  assign entriesToCheck_5_6 = _T_4766 & checkBits_5; // @[LoadQueue.scala 141:26:@4235.4]
  assign _T_4768 = storesToCheck_5_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4236.4]
  assign entriesToCheck_5_7 = _T_4768 & checkBits_5; // @[LoadQueue.scala 141:26:@4237.4]
  assign _T_4770 = storesToCheck_6_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4246.4]
  assign entriesToCheck_6_0 = _T_4770 & checkBits_6; // @[LoadQueue.scala 141:26:@4247.4]
  assign _T_4772 = storesToCheck_6_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4248.4]
  assign entriesToCheck_6_1 = _T_4772 & checkBits_6; // @[LoadQueue.scala 141:26:@4249.4]
  assign _T_4774 = storesToCheck_6_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4250.4]
  assign entriesToCheck_6_2 = _T_4774 & checkBits_6; // @[LoadQueue.scala 141:26:@4251.4]
  assign _T_4776 = storesToCheck_6_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4252.4]
  assign entriesToCheck_6_3 = _T_4776 & checkBits_6; // @[LoadQueue.scala 141:26:@4253.4]
  assign _T_4778 = storesToCheck_6_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4254.4]
  assign entriesToCheck_6_4 = _T_4778 & checkBits_6; // @[LoadQueue.scala 141:26:@4255.4]
  assign _T_4780 = storesToCheck_6_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4256.4]
  assign entriesToCheck_6_5 = _T_4780 & checkBits_6; // @[LoadQueue.scala 141:26:@4257.4]
  assign _T_4782 = storesToCheck_6_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4258.4]
  assign entriesToCheck_6_6 = _T_4782 & checkBits_6; // @[LoadQueue.scala 141:26:@4259.4]
  assign _T_4784 = storesToCheck_6_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4260.4]
  assign entriesToCheck_6_7 = _T_4784 & checkBits_6; // @[LoadQueue.scala 141:26:@4261.4]
  assign _T_4786 = storesToCheck_7_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4270.4]
  assign entriesToCheck_7_0 = _T_4786 & checkBits_7; // @[LoadQueue.scala 141:26:@4271.4]
  assign _T_4788 = storesToCheck_7_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4272.4]
  assign entriesToCheck_7_1 = _T_4788 & checkBits_7; // @[LoadQueue.scala 141:26:@4273.4]
  assign _T_4790 = storesToCheck_7_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4274.4]
  assign entriesToCheck_7_2 = _T_4790 & checkBits_7; // @[LoadQueue.scala 141:26:@4275.4]
  assign _T_4792 = storesToCheck_7_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4276.4]
  assign entriesToCheck_7_3 = _T_4792 & checkBits_7; // @[LoadQueue.scala 141:26:@4277.4]
  assign _T_4794 = storesToCheck_7_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4278.4]
  assign entriesToCheck_7_4 = _T_4794 & checkBits_7; // @[LoadQueue.scala 141:26:@4279.4]
  assign _T_4796 = storesToCheck_7_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4280.4]
  assign entriesToCheck_7_5 = _T_4796 & checkBits_7; // @[LoadQueue.scala 141:26:@4281.4]
  assign _T_4798 = storesToCheck_7_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4282.4]
  assign entriesToCheck_7_6 = _T_4798 & checkBits_7; // @[LoadQueue.scala 141:26:@4283.4]
  assign _T_4800 = storesToCheck_7_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4284.4]
  assign entriesToCheck_7_7 = _T_4800 & checkBits_7; // @[LoadQueue.scala 141:26:@4285.4]
  assign _T_5168 = entriesToCheck_0_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@4295.4]
  assign _T_5169 = _T_5168 & addrKnown_0; // @[LoadQueue.scala 152:41:@4296.4]
  assign _T_5170 = addrQ_0 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@4297.4]
  assign conflict_0_0 = _T_5169 & _T_5170; // @[LoadQueue.scala 152:68:@4298.4]
  assign _T_5172 = entriesToCheck_0_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@4300.4]
  assign _T_5173 = _T_5172 & addrKnown_0; // @[LoadQueue.scala 152:41:@4301.4]
  assign _T_5174 = addrQ_0 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@4302.4]
  assign conflict_0_1 = _T_5173 & _T_5174; // @[LoadQueue.scala 152:68:@4303.4]
  assign _T_5176 = entriesToCheck_0_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@4305.4]
  assign _T_5177 = _T_5176 & addrKnown_0; // @[LoadQueue.scala 152:41:@4306.4]
  assign _T_5178 = addrQ_0 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@4307.4]
  assign conflict_0_2 = _T_5177 & _T_5178; // @[LoadQueue.scala 152:68:@4308.4]
  assign _T_5180 = entriesToCheck_0_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@4310.4]
  assign _T_5181 = _T_5180 & addrKnown_0; // @[LoadQueue.scala 152:41:@4311.4]
  assign _T_5182 = addrQ_0 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@4312.4]
  assign conflict_0_3 = _T_5181 & _T_5182; // @[LoadQueue.scala 152:68:@4313.4]
  assign _T_5184 = entriesToCheck_0_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@4315.4]
  assign _T_5185 = _T_5184 & addrKnown_0; // @[LoadQueue.scala 152:41:@4316.4]
  assign _T_5186 = addrQ_0 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@4317.4]
  assign conflict_0_4 = _T_5185 & _T_5186; // @[LoadQueue.scala 152:68:@4318.4]
  assign _T_5188 = entriesToCheck_0_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@4320.4]
  assign _T_5189 = _T_5188 & addrKnown_0; // @[LoadQueue.scala 152:41:@4321.4]
  assign _T_5190 = addrQ_0 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@4322.4]
  assign conflict_0_5 = _T_5189 & _T_5190; // @[LoadQueue.scala 152:68:@4323.4]
  assign _T_5192 = entriesToCheck_0_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@4325.4]
  assign _T_5193 = _T_5192 & addrKnown_0; // @[LoadQueue.scala 152:41:@4326.4]
  assign _T_5194 = addrQ_0 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@4327.4]
  assign conflict_0_6 = _T_5193 & _T_5194; // @[LoadQueue.scala 152:68:@4328.4]
  assign _T_5196 = entriesToCheck_0_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@4330.4]
  assign _T_5197 = _T_5196 & addrKnown_0; // @[LoadQueue.scala 152:41:@4331.4]
  assign _T_5198 = addrQ_0 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@4332.4]
  assign conflict_0_7 = _T_5197 & _T_5198; // @[LoadQueue.scala 152:68:@4333.4]
  assign _T_5200 = entriesToCheck_1_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@4335.4]
  assign _T_5201 = _T_5200 & addrKnown_1; // @[LoadQueue.scala 152:41:@4336.4]
  assign _T_5202 = addrQ_1 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@4337.4]
  assign conflict_1_0 = _T_5201 & _T_5202; // @[LoadQueue.scala 152:68:@4338.4]
  assign _T_5204 = entriesToCheck_1_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@4340.4]
  assign _T_5205 = _T_5204 & addrKnown_1; // @[LoadQueue.scala 152:41:@4341.4]
  assign _T_5206 = addrQ_1 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@4342.4]
  assign conflict_1_1 = _T_5205 & _T_5206; // @[LoadQueue.scala 152:68:@4343.4]
  assign _T_5208 = entriesToCheck_1_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@4345.4]
  assign _T_5209 = _T_5208 & addrKnown_1; // @[LoadQueue.scala 152:41:@4346.4]
  assign _T_5210 = addrQ_1 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@4347.4]
  assign conflict_1_2 = _T_5209 & _T_5210; // @[LoadQueue.scala 152:68:@4348.4]
  assign _T_5212 = entriesToCheck_1_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@4350.4]
  assign _T_5213 = _T_5212 & addrKnown_1; // @[LoadQueue.scala 152:41:@4351.4]
  assign _T_5214 = addrQ_1 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@4352.4]
  assign conflict_1_3 = _T_5213 & _T_5214; // @[LoadQueue.scala 152:68:@4353.4]
  assign _T_5216 = entriesToCheck_1_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@4355.4]
  assign _T_5217 = _T_5216 & addrKnown_1; // @[LoadQueue.scala 152:41:@4356.4]
  assign _T_5218 = addrQ_1 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@4357.4]
  assign conflict_1_4 = _T_5217 & _T_5218; // @[LoadQueue.scala 152:68:@4358.4]
  assign _T_5220 = entriesToCheck_1_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@4360.4]
  assign _T_5221 = _T_5220 & addrKnown_1; // @[LoadQueue.scala 152:41:@4361.4]
  assign _T_5222 = addrQ_1 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@4362.4]
  assign conflict_1_5 = _T_5221 & _T_5222; // @[LoadQueue.scala 152:68:@4363.4]
  assign _T_5224 = entriesToCheck_1_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@4365.4]
  assign _T_5225 = _T_5224 & addrKnown_1; // @[LoadQueue.scala 152:41:@4366.4]
  assign _T_5226 = addrQ_1 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@4367.4]
  assign conflict_1_6 = _T_5225 & _T_5226; // @[LoadQueue.scala 152:68:@4368.4]
  assign _T_5228 = entriesToCheck_1_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@4370.4]
  assign _T_5229 = _T_5228 & addrKnown_1; // @[LoadQueue.scala 152:41:@4371.4]
  assign _T_5230 = addrQ_1 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@4372.4]
  assign conflict_1_7 = _T_5229 & _T_5230; // @[LoadQueue.scala 152:68:@4373.4]
  assign _T_5232 = entriesToCheck_2_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@4375.4]
  assign _T_5233 = _T_5232 & addrKnown_2; // @[LoadQueue.scala 152:41:@4376.4]
  assign _T_5234 = addrQ_2 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@4377.4]
  assign conflict_2_0 = _T_5233 & _T_5234; // @[LoadQueue.scala 152:68:@4378.4]
  assign _T_5236 = entriesToCheck_2_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@4380.4]
  assign _T_5237 = _T_5236 & addrKnown_2; // @[LoadQueue.scala 152:41:@4381.4]
  assign _T_5238 = addrQ_2 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@4382.4]
  assign conflict_2_1 = _T_5237 & _T_5238; // @[LoadQueue.scala 152:68:@4383.4]
  assign _T_5240 = entriesToCheck_2_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@4385.4]
  assign _T_5241 = _T_5240 & addrKnown_2; // @[LoadQueue.scala 152:41:@4386.4]
  assign _T_5242 = addrQ_2 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@4387.4]
  assign conflict_2_2 = _T_5241 & _T_5242; // @[LoadQueue.scala 152:68:@4388.4]
  assign _T_5244 = entriesToCheck_2_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@4390.4]
  assign _T_5245 = _T_5244 & addrKnown_2; // @[LoadQueue.scala 152:41:@4391.4]
  assign _T_5246 = addrQ_2 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@4392.4]
  assign conflict_2_3 = _T_5245 & _T_5246; // @[LoadQueue.scala 152:68:@4393.4]
  assign _T_5248 = entriesToCheck_2_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@4395.4]
  assign _T_5249 = _T_5248 & addrKnown_2; // @[LoadQueue.scala 152:41:@4396.4]
  assign _T_5250 = addrQ_2 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@4397.4]
  assign conflict_2_4 = _T_5249 & _T_5250; // @[LoadQueue.scala 152:68:@4398.4]
  assign _T_5252 = entriesToCheck_2_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@4400.4]
  assign _T_5253 = _T_5252 & addrKnown_2; // @[LoadQueue.scala 152:41:@4401.4]
  assign _T_5254 = addrQ_2 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@4402.4]
  assign conflict_2_5 = _T_5253 & _T_5254; // @[LoadQueue.scala 152:68:@4403.4]
  assign _T_5256 = entriesToCheck_2_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@4405.4]
  assign _T_5257 = _T_5256 & addrKnown_2; // @[LoadQueue.scala 152:41:@4406.4]
  assign _T_5258 = addrQ_2 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@4407.4]
  assign conflict_2_6 = _T_5257 & _T_5258; // @[LoadQueue.scala 152:68:@4408.4]
  assign _T_5260 = entriesToCheck_2_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@4410.4]
  assign _T_5261 = _T_5260 & addrKnown_2; // @[LoadQueue.scala 152:41:@4411.4]
  assign _T_5262 = addrQ_2 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@4412.4]
  assign conflict_2_7 = _T_5261 & _T_5262; // @[LoadQueue.scala 152:68:@4413.4]
  assign _T_5264 = entriesToCheck_3_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@4415.4]
  assign _T_5265 = _T_5264 & addrKnown_3; // @[LoadQueue.scala 152:41:@4416.4]
  assign _T_5266 = addrQ_3 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@4417.4]
  assign conflict_3_0 = _T_5265 & _T_5266; // @[LoadQueue.scala 152:68:@4418.4]
  assign _T_5268 = entriesToCheck_3_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@4420.4]
  assign _T_5269 = _T_5268 & addrKnown_3; // @[LoadQueue.scala 152:41:@4421.4]
  assign _T_5270 = addrQ_3 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@4422.4]
  assign conflict_3_1 = _T_5269 & _T_5270; // @[LoadQueue.scala 152:68:@4423.4]
  assign _T_5272 = entriesToCheck_3_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@4425.4]
  assign _T_5273 = _T_5272 & addrKnown_3; // @[LoadQueue.scala 152:41:@4426.4]
  assign _T_5274 = addrQ_3 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@4427.4]
  assign conflict_3_2 = _T_5273 & _T_5274; // @[LoadQueue.scala 152:68:@4428.4]
  assign _T_5276 = entriesToCheck_3_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@4430.4]
  assign _T_5277 = _T_5276 & addrKnown_3; // @[LoadQueue.scala 152:41:@4431.4]
  assign _T_5278 = addrQ_3 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@4432.4]
  assign conflict_3_3 = _T_5277 & _T_5278; // @[LoadQueue.scala 152:68:@4433.4]
  assign _T_5280 = entriesToCheck_3_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@4435.4]
  assign _T_5281 = _T_5280 & addrKnown_3; // @[LoadQueue.scala 152:41:@4436.4]
  assign _T_5282 = addrQ_3 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@4437.4]
  assign conflict_3_4 = _T_5281 & _T_5282; // @[LoadQueue.scala 152:68:@4438.4]
  assign _T_5284 = entriesToCheck_3_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@4440.4]
  assign _T_5285 = _T_5284 & addrKnown_3; // @[LoadQueue.scala 152:41:@4441.4]
  assign _T_5286 = addrQ_3 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@4442.4]
  assign conflict_3_5 = _T_5285 & _T_5286; // @[LoadQueue.scala 152:68:@4443.4]
  assign _T_5288 = entriesToCheck_3_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@4445.4]
  assign _T_5289 = _T_5288 & addrKnown_3; // @[LoadQueue.scala 152:41:@4446.4]
  assign _T_5290 = addrQ_3 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@4447.4]
  assign conflict_3_6 = _T_5289 & _T_5290; // @[LoadQueue.scala 152:68:@4448.4]
  assign _T_5292 = entriesToCheck_3_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@4450.4]
  assign _T_5293 = _T_5292 & addrKnown_3; // @[LoadQueue.scala 152:41:@4451.4]
  assign _T_5294 = addrQ_3 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@4452.4]
  assign conflict_3_7 = _T_5293 & _T_5294; // @[LoadQueue.scala 152:68:@4453.4]
  assign _T_5296 = entriesToCheck_4_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@4455.4]
  assign _T_5297 = _T_5296 & addrKnown_4; // @[LoadQueue.scala 152:41:@4456.4]
  assign _T_5298 = addrQ_4 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@4457.4]
  assign conflict_4_0 = _T_5297 & _T_5298; // @[LoadQueue.scala 152:68:@4458.4]
  assign _T_5300 = entriesToCheck_4_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@4460.4]
  assign _T_5301 = _T_5300 & addrKnown_4; // @[LoadQueue.scala 152:41:@4461.4]
  assign _T_5302 = addrQ_4 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@4462.4]
  assign conflict_4_1 = _T_5301 & _T_5302; // @[LoadQueue.scala 152:68:@4463.4]
  assign _T_5304 = entriesToCheck_4_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@4465.4]
  assign _T_5305 = _T_5304 & addrKnown_4; // @[LoadQueue.scala 152:41:@4466.4]
  assign _T_5306 = addrQ_4 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@4467.4]
  assign conflict_4_2 = _T_5305 & _T_5306; // @[LoadQueue.scala 152:68:@4468.4]
  assign _T_5308 = entriesToCheck_4_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@4470.4]
  assign _T_5309 = _T_5308 & addrKnown_4; // @[LoadQueue.scala 152:41:@4471.4]
  assign _T_5310 = addrQ_4 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@4472.4]
  assign conflict_4_3 = _T_5309 & _T_5310; // @[LoadQueue.scala 152:68:@4473.4]
  assign _T_5312 = entriesToCheck_4_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@4475.4]
  assign _T_5313 = _T_5312 & addrKnown_4; // @[LoadQueue.scala 152:41:@4476.4]
  assign _T_5314 = addrQ_4 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@4477.4]
  assign conflict_4_4 = _T_5313 & _T_5314; // @[LoadQueue.scala 152:68:@4478.4]
  assign _T_5316 = entriesToCheck_4_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@4480.4]
  assign _T_5317 = _T_5316 & addrKnown_4; // @[LoadQueue.scala 152:41:@4481.4]
  assign _T_5318 = addrQ_4 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@4482.4]
  assign conflict_4_5 = _T_5317 & _T_5318; // @[LoadQueue.scala 152:68:@4483.4]
  assign _T_5320 = entriesToCheck_4_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@4485.4]
  assign _T_5321 = _T_5320 & addrKnown_4; // @[LoadQueue.scala 152:41:@4486.4]
  assign _T_5322 = addrQ_4 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@4487.4]
  assign conflict_4_6 = _T_5321 & _T_5322; // @[LoadQueue.scala 152:68:@4488.4]
  assign _T_5324 = entriesToCheck_4_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@4490.4]
  assign _T_5325 = _T_5324 & addrKnown_4; // @[LoadQueue.scala 152:41:@4491.4]
  assign _T_5326 = addrQ_4 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@4492.4]
  assign conflict_4_7 = _T_5325 & _T_5326; // @[LoadQueue.scala 152:68:@4493.4]
  assign _T_5328 = entriesToCheck_5_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@4495.4]
  assign _T_5329 = _T_5328 & addrKnown_5; // @[LoadQueue.scala 152:41:@4496.4]
  assign _T_5330 = addrQ_5 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@4497.4]
  assign conflict_5_0 = _T_5329 & _T_5330; // @[LoadQueue.scala 152:68:@4498.4]
  assign _T_5332 = entriesToCheck_5_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@4500.4]
  assign _T_5333 = _T_5332 & addrKnown_5; // @[LoadQueue.scala 152:41:@4501.4]
  assign _T_5334 = addrQ_5 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@4502.4]
  assign conflict_5_1 = _T_5333 & _T_5334; // @[LoadQueue.scala 152:68:@4503.4]
  assign _T_5336 = entriesToCheck_5_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@4505.4]
  assign _T_5337 = _T_5336 & addrKnown_5; // @[LoadQueue.scala 152:41:@4506.4]
  assign _T_5338 = addrQ_5 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@4507.4]
  assign conflict_5_2 = _T_5337 & _T_5338; // @[LoadQueue.scala 152:68:@4508.4]
  assign _T_5340 = entriesToCheck_5_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@4510.4]
  assign _T_5341 = _T_5340 & addrKnown_5; // @[LoadQueue.scala 152:41:@4511.4]
  assign _T_5342 = addrQ_5 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@4512.4]
  assign conflict_5_3 = _T_5341 & _T_5342; // @[LoadQueue.scala 152:68:@4513.4]
  assign _T_5344 = entriesToCheck_5_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@4515.4]
  assign _T_5345 = _T_5344 & addrKnown_5; // @[LoadQueue.scala 152:41:@4516.4]
  assign _T_5346 = addrQ_5 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@4517.4]
  assign conflict_5_4 = _T_5345 & _T_5346; // @[LoadQueue.scala 152:68:@4518.4]
  assign _T_5348 = entriesToCheck_5_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@4520.4]
  assign _T_5349 = _T_5348 & addrKnown_5; // @[LoadQueue.scala 152:41:@4521.4]
  assign _T_5350 = addrQ_5 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@4522.4]
  assign conflict_5_5 = _T_5349 & _T_5350; // @[LoadQueue.scala 152:68:@4523.4]
  assign _T_5352 = entriesToCheck_5_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@4525.4]
  assign _T_5353 = _T_5352 & addrKnown_5; // @[LoadQueue.scala 152:41:@4526.4]
  assign _T_5354 = addrQ_5 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@4527.4]
  assign conflict_5_6 = _T_5353 & _T_5354; // @[LoadQueue.scala 152:68:@4528.4]
  assign _T_5356 = entriesToCheck_5_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@4530.4]
  assign _T_5357 = _T_5356 & addrKnown_5; // @[LoadQueue.scala 152:41:@4531.4]
  assign _T_5358 = addrQ_5 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@4532.4]
  assign conflict_5_7 = _T_5357 & _T_5358; // @[LoadQueue.scala 152:68:@4533.4]
  assign _T_5360 = entriesToCheck_6_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@4535.4]
  assign _T_5361 = _T_5360 & addrKnown_6; // @[LoadQueue.scala 152:41:@4536.4]
  assign _T_5362 = addrQ_6 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@4537.4]
  assign conflict_6_0 = _T_5361 & _T_5362; // @[LoadQueue.scala 152:68:@4538.4]
  assign _T_5364 = entriesToCheck_6_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@4540.4]
  assign _T_5365 = _T_5364 & addrKnown_6; // @[LoadQueue.scala 152:41:@4541.4]
  assign _T_5366 = addrQ_6 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@4542.4]
  assign conflict_6_1 = _T_5365 & _T_5366; // @[LoadQueue.scala 152:68:@4543.4]
  assign _T_5368 = entriesToCheck_6_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@4545.4]
  assign _T_5369 = _T_5368 & addrKnown_6; // @[LoadQueue.scala 152:41:@4546.4]
  assign _T_5370 = addrQ_6 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@4547.4]
  assign conflict_6_2 = _T_5369 & _T_5370; // @[LoadQueue.scala 152:68:@4548.4]
  assign _T_5372 = entriesToCheck_6_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@4550.4]
  assign _T_5373 = _T_5372 & addrKnown_6; // @[LoadQueue.scala 152:41:@4551.4]
  assign _T_5374 = addrQ_6 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@4552.4]
  assign conflict_6_3 = _T_5373 & _T_5374; // @[LoadQueue.scala 152:68:@4553.4]
  assign _T_5376 = entriesToCheck_6_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@4555.4]
  assign _T_5377 = _T_5376 & addrKnown_6; // @[LoadQueue.scala 152:41:@4556.4]
  assign _T_5378 = addrQ_6 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@4557.4]
  assign conflict_6_4 = _T_5377 & _T_5378; // @[LoadQueue.scala 152:68:@4558.4]
  assign _T_5380 = entriesToCheck_6_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@4560.4]
  assign _T_5381 = _T_5380 & addrKnown_6; // @[LoadQueue.scala 152:41:@4561.4]
  assign _T_5382 = addrQ_6 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@4562.4]
  assign conflict_6_5 = _T_5381 & _T_5382; // @[LoadQueue.scala 152:68:@4563.4]
  assign _T_5384 = entriesToCheck_6_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@4565.4]
  assign _T_5385 = _T_5384 & addrKnown_6; // @[LoadQueue.scala 152:41:@4566.4]
  assign _T_5386 = addrQ_6 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@4567.4]
  assign conflict_6_6 = _T_5385 & _T_5386; // @[LoadQueue.scala 152:68:@4568.4]
  assign _T_5388 = entriesToCheck_6_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@4570.4]
  assign _T_5389 = _T_5388 & addrKnown_6; // @[LoadQueue.scala 152:41:@4571.4]
  assign _T_5390 = addrQ_6 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@4572.4]
  assign conflict_6_7 = _T_5389 & _T_5390; // @[LoadQueue.scala 152:68:@4573.4]
  assign _T_5392 = entriesToCheck_7_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@4575.4]
  assign _T_5393 = _T_5392 & addrKnown_7; // @[LoadQueue.scala 152:41:@4576.4]
  assign _T_5394 = addrQ_7 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@4577.4]
  assign conflict_7_0 = _T_5393 & _T_5394; // @[LoadQueue.scala 152:68:@4578.4]
  assign _T_5396 = entriesToCheck_7_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@4580.4]
  assign _T_5397 = _T_5396 & addrKnown_7; // @[LoadQueue.scala 152:41:@4581.4]
  assign _T_5398 = addrQ_7 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@4582.4]
  assign conflict_7_1 = _T_5397 & _T_5398; // @[LoadQueue.scala 152:68:@4583.4]
  assign _T_5400 = entriesToCheck_7_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@4585.4]
  assign _T_5401 = _T_5400 & addrKnown_7; // @[LoadQueue.scala 152:41:@4586.4]
  assign _T_5402 = addrQ_7 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@4587.4]
  assign conflict_7_2 = _T_5401 & _T_5402; // @[LoadQueue.scala 152:68:@4588.4]
  assign _T_5404 = entriesToCheck_7_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@4590.4]
  assign _T_5405 = _T_5404 & addrKnown_7; // @[LoadQueue.scala 152:41:@4591.4]
  assign _T_5406 = addrQ_7 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@4592.4]
  assign conflict_7_3 = _T_5405 & _T_5406; // @[LoadQueue.scala 152:68:@4593.4]
  assign _T_5408 = entriesToCheck_7_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@4595.4]
  assign _T_5409 = _T_5408 & addrKnown_7; // @[LoadQueue.scala 152:41:@4596.4]
  assign _T_5410 = addrQ_7 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@4597.4]
  assign conflict_7_4 = _T_5409 & _T_5410; // @[LoadQueue.scala 152:68:@4598.4]
  assign _T_5412 = entriesToCheck_7_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@4600.4]
  assign _T_5413 = _T_5412 & addrKnown_7; // @[LoadQueue.scala 152:41:@4601.4]
  assign _T_5414 = addrQ_7 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@4602.4]
  assign conflict_7_5 = _T_5413 & _T_5414; // @[LoadQueue.scala 152:68:@4603.4]
  assign _T_5416 = entriesToCheck_7_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@4605.4]
  assign _T_5417 = _T_5416 & addrKnown_7; // @[LoadQueue.scala 152:41:@4606.4]
  assign _T_5418 = addrQ_7 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@4607.4]
  assign conflict_7_6 = _T_5417 & _T_5418; // @[LoadQueue.scala 152:68:@4608.4]
  assign _T_5420 = entriesToCheck_7_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@4610.4]
  assign _T_5421 = _T_5420 & addrKnown_7; // @[LoadQueue.scala 152:41:@4611.4]
  assign _T_5422 = addrQ_7 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@4612.4]
  assign conflict_7_7 = _T_5421 & _T_5422; // @[LoadQueue.scala 152:68:@4613.4]
  assign _T_5791 = io_storeAddrDone_0 == 1'h0; // @[LoadQueue.scala 163:13:@4616.4]
  assign storeAddrNotKnownFlags_0_0 = _T_5791 & entriesToCheck_0_0; // @[LoadQueue.scala 163:19:@4617.4]
  assign _T_5794 = io_storeAddrDone_1 == 1'h0; // @[LoadQueue.scala 163:13:@4618.4]
  assign storeAddrNotKnownFlags_0_1 = _T_5794 & entriesToCheck_0_1; // @[LoadQueue.scala 163:19:@4619.4]
  assign _T_5797 = io_storeAddrDone_2 == 1'h0; // @[LoadQueue.scala 163:13:@4620.4]
  assign storeAddrNotKnownFlags_0_2 = _T_5797 & entriesToCheck_0_2; // @[LoadQueue.scala 163:19:@4621.4]
  assign _T_5800 = io_storeAddrDone_3 == 1'h0; // @[LoadQueue.scala 163:13:@4622.4]
  assign storeAddrNotKnownFlags_0_3 = _T_5800 & entriesToCheck_0_3; // @[LoadQueue.scala 163:19:@4623.4]
  assign _T_5803 = io_storeAddrDone_4 == 1'h0; // @[LoadQueue.scala 163:13:@4624.4]
  assign storeAddrNotKnownFlags_0_4 = _T_5803 & entriesToCheck_0_4; // @[LoadQueue.scala 163:19:@4625.4]
  assign _T_5806 = io_storeAddrDone_5 == 1'h0; // @[LoadQueue.scala 163:13:@4626.4]
  assign storeAddrNotKnownFlags_0_5 = _T_5806 & entriesToCheck_0_5; // @[LoadQueue.scala 163:19:@4627.4]
  assign _T_5809 = io_storeAddrDone_6 == 1'h0; // @[LoadQueue.scala 163:13:@4628.4]
  assign storeAddrNotKnownFlags_0_6 = _T_5809 & entriesToCheck_0_6; // @[LoadQueue.scala 163:19:@4629.4]
  assign _T_5812 = io_storeAddrDone_7 == 1'h0; // @[LoadQueue.scala 163:13:@4630.4]
  assign storeAddrNotKnownFlags_0_7 = _T_5812 & entriesToCheck_0_7; // @[LoadQueue.scala 163:19:@4631.4]
  assign storeAddrNotKnownFlags_1_0 = _T_5791 & entriesToCheck_1_0; // @[LoadQueue.scala 163:19:@4641.4]
  assign storeAddrNotKnownFlags_1_1 = _T_5794 & entriesToCheck_1_1; // @[LoadQueue.scala 163:19:@4643.4]
  assign storeAddrNotKnownFlags_1_2 = _T_5797 & entriesToCheck_1_2; // @[LoadQueue.scala 163:19:@4645.4]
  assign storeAddrNotKnownFlags_1_3 = _T_5800 & entriesToCheck_1_3; // @[LoadQueue.scala 163:19:@4647.4]
  assign storeAddrNotKnownFlags_1_4 = _T_5803 & entriesToCheck_1_4; // @[LoadQueue.scala 163:19:@4649.4]
  assign storeAddrNotKnownFlags_1_5 = _T_5806 & entriesToCheck_1_5; // @[LoadQueue.scala 163:19:@4651.4]
  assign storeAddrNotKnownFlags_1_6 = _T_5809 & entriesToCheck_1_6; // @[LoadQueue.scala 163:19:@4653.4]
  assign storeAddrNotKnownFlags_1_7 = _T_5812 & entriesToCheck_1_7; // @[LoadQueue.scala 163:19:@4655.4]
  assign storeAddrNotKnownFlags_2_0 = _T_5791 & entriesToCheck_2_0; // @[LoadQueue.scala 163:19:@4665.4]
  assign storeAddrNotKnownFlags_2_1 = _T_5794 & entriesToCheck_2_1; // @[LoadQueue.scala 163:19:@4667.4]
  assign storeAddrNotKnownFlags_2_2 = _T_5797 & entriesToCheck_2_2; // @[LoadQueue.scala 163:19:@4669.4]
  assign storeAddrNotKnownFlags_2_3 = _T_5800 & entriesToCheck_2_3; // @[LoadQueue.scala 163:19:@4671.4]
  assign storeAddrNotKnownFlags_2_4 = _T_5803 & entriesToCheck_2_4; // @[LoadQueue.scala 163:19:@4673.4]
  assign storeAddrNotKnownFlags_2_5 = _T_5806 & entriesToCheck_2_5; // @[LoadQueue.scala 163:19:@4675.4]
  assign storeAddrNotKnownFlags_2_6 = _T_5809 & entriesToCheck_2_6; // @[LoadQueue.scala 163:19:@4677.4]
  assign storeAddrNotKnownFlags_2_7 = _T_5812 & entriesToCheck_2_7; // @[LoadQueue.scala 163:19:@4679.4]
  assign storeAddrNotKnownFlags_3_0 = _T_5791 & entriesToCheck_3_0; // @[LoadQueue.scala 163:19:@4689.4]
  assign storeAddrNotKnownFlags_3_1 = _T_5794 & entriesToCheck_3_1; // @[LoadQueue.scala 163:19:@4691.4]
  assign storeAddrNotKnownFlags_3_2 = _T_5797 & entriesToCheck_3_2; // @[LoadQueue.scala 163:19:@4693.4]
  assign storeAddrNotKnownFlags_3_3 = _T_5800 & entriesToCheck_3_3; // @[LoadQueue.scala 163:19:@4695.4]
  assign storeAddrNotKnownFlags_3_4 = _T_5803 & entriesToCheck_3_4; // @[LoadQueue.scala 163:19:@4697.4]
  assign storeAddrNotKnownFlags_3_5 = _T_5806 & entriesToCheck_3_5; // @[LoadQueue.scala 163:19:@4699.4]
  assign storeAddrNotKnownFlags_3_6 = _T_5809 & entriesToCheck_3_6; // @[LoadQueue.scala 163:19:@4701.4]
  assign storeAddrNotKnownFlags_3_7 = _T_5812 & entriesToCheck_3_7; // @[LoadQueue.scala 163:19:@4703.4]
  assign storeAddrNotKnownFlags_4_0 = _T_5791 & entriesToCheck_4_0; // @[LoadQueue.scala 163:19:@4713.4]
  assign storeAddrNotKnownFlags_4_1 = _T_5794 & entriesToCheck_4_1; // @[LoadQueue.scala 163:19:@4715.4]
  assign storeAddrNotKnownFlags_4_2 = _T_5797 & entriesToCheck_4_2; // @[LoadQueue.scala 163:19:@4717.4]
  assign storeAddrNotKnownFlags_4_3 = _T_5800 & entriesToCheck_4_3; // @[LoadQueue.scala 163:19:@4719.4]
  assign storeAddrNotKnownFlags_4_4 = _T_5803 & entriesToCheck_4_4; // @[LoadQueue.scala 163:19:@4721.4]
  assign storeAddrNotKnownFlags_4_5 = _T_5806 & entriesToCheck_4_5; // @[LoadQueue.scala 163:19:@4723.4]
  assign storeAddrNotKnownFlags_4_6 = _T_5809 & entriesToCheck_4_6; // @[LoadQueue.scala 163:19:@4725.4]
  assign storeAddrNotKnownFlags_4_7 = _T_5812 & entriesToCheck_4_7; // @[LoadQueue.scala 163:19:@4727.4]
  assign storeAddrNotKnownFlags_5_0 = _T_5791 & entriesToCheck_5_0; // @[LoadQueue.scala 163:19:@4737.4]
  assign storeAddrNotKnownFlags_5_1 = _T_5794 & entriesToCheck_5_1; // @[LoadQueue.scala 163:19:@4739.4]
  assign storeAddrNotKnownFlags_5_2 = _T_5797 & entriesToCheck_5_2; // @[LoadQueue.scala 163:19:@4741.4]
  assign storeAddrNotKnownFlags_5_3 = _T_5800 & entriesToCheck_5_3; // @[LoadQueue.scala 163:19:@4743.4]
  assign storeAddrNotKnownFlags_5_4 = _T_5803 & entriesToCheck_5_4; // @[LoadQueue.scala 163:19:@4745.4]
  assign storeAddrNotKnownFlags_5_5 = _T_5806 & entriesToCheck_5_5; // @[LoadQueue.scala 163:19:@4747.4]
  assign storeAddrNotKnownFlags_5_6 = _T_5809 & entriesToCheck_5_6; // @[LoadQueue.scala 163:19:@4749.4]
  assign storeAddrNotKnownFlags_5_7 = _T_5812 & entriesToCheck_5_7; // @[LoadQueue.scala 163:19:@4751.4]
  assign storeAddrNotKnownFlags_6_0 = _T_5791 & entriesToCheck_6_0; // @[LoadQueue.scala 163:19:@4761.4]
  assign storeAddrNotKnownFlags_6_1 = _T_5794 & entriesToCheck_6_1; // @[LoadQueue.scala 163:19:@4763.4]
  assign storeAddrNotKnownFlags_6_2 = _T_5797 & entriesToCheck_6_2; // @[LoadQueue.scala 163:19:@4765.4]
  assign storeAddrNotKnownFlags_6_3 = _T_5800 & entriesToCheck_6_3; // @[LoadQueue.scala 163:19:@4767.4]
  assign storeAddrNotKnownFlags_6_4 = _T_5803 & entriesToCheck_6_4; // @[LoadQueue.scala 163:19:@4769.4]
  assign storeAddrNotKnownFlags_6_5 = _T_5806 & entriesToCheck_6_5; // @[LoadQueue.scala 163:19:@4771.4]
  assign storeAddrNotKnownFlags_6_6 = _T_5809 & entriesToCheck_6_6; // @[LoadQueue.scala 163:19:@4773.4]
  assign storeAddrNotKnownFlags_6_7 = _T_5812 & entriesToCheck_6_7; // @[LoadQueue.scala 163:19:@4775.4]
  assign storeAddrNotKnownFlags_7_0 = _T_5791 & entriesToCheck_7_0; // @[LoadQueue.scala 163:19:@4785.4]
  assign storeAddrNotKnownFlags_7_1 = _T_5794 & entriesToCheck_7_1; // @[LoadQueue.scala 163:19:@4787.4]
  assign storeAddrNotKnownFlags_7_2 = _T_5797 & entriesToCheck_7_2; // @[LoadQueue.scala 163:19:@4789.4]
  assign storeAddrNotKnownFlags_7_3 = _T_5800 & entriesToCheck_7_3; // @[LoadQueue.scala 163:19:@4791.4]
  assign storeAddrNotKnownFlags_7_4 = _T_5803 & entriesToCheck_7_4; // @[LoadQueue.scala 163:19:@4793.4]
  assign storeAddrNotKnownFlags_7_5 = _T_5806 & entriesToCheck_7_5; // @[LoadQueue.scala 163:19:@4795.4]
  assign storeAddrNotKnownFlags_7_6 = _T_5809 & entriesToCheck_7_6; // @[LoadQueue.scala 163:19:@4797.4]
  assign storeAddrNotKnownFlags_7_7 = _T_5812 & entriesToCheck_7_7; // @[LoadQueue.scala 163:19:@4799.4]
  assign _T_6146 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0}; // @[Mux.scala 19:72:@4906.4]
  assign _T_6148 = _T_1537 ? _T_6146 : 8'h0; // @[Mux.scala 19:72:@4907.4]
  assign _T_6155 = {conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1}; // @[Mux.scala 19:72:@4914.4]
  assign _T_6157 = _T_1538 ? _T_6155 : 8'h0; // @[Mux.scala 19:72:@4915.4]
  assign _T_6164 = {conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2}; // @[Mux.scala 19:72:@4922.4]
  assign _T_6166 = _T_1539 ? _T_6164 : 8'h0; // @[Mux.scala 19:72:@4923.4]
  assign _T_6173 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3}; // @[Mux.scala 19:72:@4930.4]
  assign _T_6175 = _T_1540 ? _T_6173 : 8'h0; // @[Mux.scala 19:72:@4931.4]
  assign _T_6182 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4}; // @[Mux.scala 19:72:@4938.4]
  assign _T_6184 = _T_1541 ? _T_6182 : 8'h0; // @[Mux.scala 19:72:@4939.4]
  assign _T_6191 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5}; // @[Mux.scala 19:72:@4946.4]
  assign _T_6193 = _T_1542 ? _T_6191 : 8'h0; // @[Mux.scala 19:72:@4947.4]
  assign _T_6200 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6}; // @[Mux.scala 19:72:@4954.4]
  assign _T_6202 = _T_1543 ? _T_6200 : 8'h0; // @[Mux.scala 19:72:@4955.4]
  assign _T_6209 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7}; // @[Mux.scala 19:72:@4962.4]
  assign _T_6211 = _T_1544 ? _T_6209 : 8'h0; // @[Mux.scala 19:72:@4963.4]
  assign _T_6212 = _T_6148 | _T_6157; // @[Mux.scala 19:72:@4964.4]
  assign _T_6213 = _T_6212 | _T_6166; // @[Mux.scala 19:72:@4965.4]
  assign _T_6214 = _T_6213 | _T_6175; // @[Mux.scala 19:72:@4966.4]
  assign _T_6215 = _T_6214 | _T_6184; // @[Mux.scala 19:72:@4967.4]
  assign _T_6216 = _T_6215 | _T_6193; // @[Mux.scala 19:72:@4968.4]
  assign _T_6217 = _T_6216 | _T_6202; // @[Mux.scala 19:72:@4969.4]
  assign _T_6218 = _T_6217 | _T_6211; // @[Mux.scala 19:72:@4970.4]
  assign _T_6460 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0}; // @[Mux.scala 19:72:@5088.4]
  assign _T_6462 = _T_1537 ? _T_6460 : 8'h0; // @[Mux.scala 19:72:@5089.4]
  assign _T_6469 = {conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1}; // @[Mux.scala 19:72:@5096.4]
  assign _T_6471 = _T_1538 ? _T_6469 : 8'h0; // @[Mux.scala 19:72:@5097.4]
  assign _T_6478 = {conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2}; // @[Mux.scala 19:72:@5104.4]
  assign _T_6480 = _T_1539 ? _T_6478 : 8'h0; // @[Mux.scala 19:72:@5105.4]
  assign _T_6487 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3}; // @[Mux.scala 19:72:@5112.4]
  assign _T_6489 = _T_1540 ? _T_6487 : 8'h0; // @[Mux.scala 19:72:@5113.4]
  assign _T_6496 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4}; // @[Mux.scala 19:72:@5120.4]
  assign _T_6498 = _T_1541 ? _T_6496 : 8'h0; // @[Mux.scala 19:72:@5121.4]
  assign _T_6505 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5}; // @[Mux.scala 19:72:@5128.4]
  assign _T_6507 = _T_1542 ? _T_6505 : 8'h0; // @[Mux.scala 19:72:@5129.4]
  assign _T_6514 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6}; // @[Mux.scala 19:72:@5136.4]
  assign _T_6516 = _T_1543 ? _T_6514 : 8'h0; // @[Mux.scala 19:72:@5137.4]
  assign _T_6523 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7}; // @[Mux.scala 19:72:@5144.4]
  assign _T_6525 = _T_1544 ? _T_6523 : 8'h0; // @[Mux.scala 19:72:@5145.4]
  assign _T_6526 = _T_6462 | _T_6471; // @[Mux.scala 19:72:@5146.4]
  assign _T_6527 = _T_6526 | _T_6480; // @[Mux.scala 19:72:@5147.4]
  assign _T_6528 = _T_6527 | _T_6489; // @[Mux.scala 19:72:@5148.4]
  assign _T_6529 = _T_6528 | _T_6498; // @[Mux.scala 19:72:@5149.4]
  assign _T_6530 = _T_6529 | _T_6507; // @[Mux.scala 19:72:@5150.4]
  assign _T_6531 = _T_6530 | _T_6516; // @[Mux.scala 19:72:@5151.4]
  assign _T_6532 = _T_6531 | _T_6525; // @[Mux.scala 19:72:@5152.4]
  assign _T_6774 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0}; // @[Mux.scala 19:72:@5270.4]
  assign _T_6776 = _T_1537 ? _T_6774 : 8'h0; // @[Mux.scala 19:72:@5271.4]
  assign _T_6783 = {conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1}; // @[Mux.scala 19:72:@5278.4]
  assign _T_6785 = _T_1538 ? _T_6783 : 8'h0; // @[Mux.scala 19:72:@5279.4]
  assign _T_6792 = {conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2}; // @[Mux.scala 19:72:@5286.4]
  assign _T_6794 = _T_1539 ? _T_6792 : 8'h0; // @[Mux.scala 19:72:@5287.4]
  assign _T_6801 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3}; // @[Mux.scala 19:72:@5294.4]
  assign _T_6803 = _T_1540 ? _T_6801 : 8'h0; // @[Mux.scala 19:72:@5295.4]
  assign _T_6810 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4}; // @[Mux.scala 19:72:@5302.4]
  assign _T_6812 = _T_1541 ? _T_6810 : 8'h0; // @[Mux.scala 19:72:@5303.4]
  assign _T_6819 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5}; // @[Mux.scala 19:72:@5310.4]
  assign _T_6821 = _T_1542 ? _T_6819 : 8'h0; // @[Mux.scala 19:72:@5311.4]
  assign _T_6828 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6}; // @[Mux.scala 19:72:@5318.4]
  assign _T_6830 = _T_1543 ? _T_6828 : 8'h0; // @[Mux.scala 19:72:@5319.4]
  assign _T_6837 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7}; // @[Mux.scala 19:72:@5326.4]
  assign _T_6839 = _T_1544 ? _T_6837 : 8'h0; // @[Mux.scala 19:72:@5327.4]
  assign _T_6840 = _T_6776 | _T_6785; // @[Mux.scala 19:72:@5328.4]
  assign _T_6841 = _T_6840 | _T_6794; // @[Mux.scala 19:72:@5329.4]
  assign _T_6842 = _T_6841 | _T_6803; // @[Mux.scala 19:72:@5330.4]
  assign _T_6843 = _T_6842 | _T_6812; // @[Mux.scala 19:72:@5331.4]
  assign _T_6844 = _T_6843 | _T_6821; // @[Mux.scala 19:72:@5332.4]
  assign _T_6845 = _T_6844 | _T_6830; // @[Mux.scala 19:72:@5333.4]
  assign _T_6846 = _T_6845 | _T_6839; // @[Mux.scala 19:72:@5334.4]
  assign _T_7088 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0}; // @[Mux.scala 19:72:@5452.4]
  assign _T_7090 = _T_1537 ? _T_7088 : 8'h0; // @[Mux.scala 19:72:@5453.4]
  assign _T_7097 = {conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1}; // @[Mux.scala 19:72:@5460.4]
  assign _T_7099 = _T_1538 ? _T_7097 : 8'h0; // @[Mux.scala 19:72:@5461.4]
  assign _T_7106 = {conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2}; // @[Mux.scala 19:72:@5468.4]
  assign _T_7108 = _T_1539 ? _T_7106 : 8'h0; // @[Mux.scala 19:72:@5469.4]
  assign _T_7115 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3}; // @[Mux.scala 19:72:@5476.4]
  assign _T_7117 = _T_1540 ? _T_7115 : 8'h0; // @[Mux.scala 19:72:@5477.4]
  assign _T_7124 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4}; // @[Mux.scala 19:72:@5484.4]
  assign _T_7126 = _T_1541 ? _T_7124 : 8'h0; // @[Mux.scala 19:72:@5485.4]
  assign _T_7133 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5}; // @[Mux.scala 19:72:@5492.4]
  assign _T_7135 = _T_1542 ? _T_7133 : 8'h0; // @[Mux.scala 19:72:@5493.4]
  assign _T_7142 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6}; // @[Mux.scala 19:72:@5500.4]
  assign _T_7144 = _T_1543 ? _T_7142 : 8'h0; // @[Mux.scala 19:72:@5501.4]
  assign _T_7151 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7}; // @[Mux.scala 19:72:@5508.4]
  assign _T_7153 = _T_1544 ? _T_7151 : 8'h0; // @[Mux.scala 19:72:@5509.4]
  assign _T_7154 = _T_7090 | _T_7099; // @[Mux.scala 19:72:@5510.4]
  assign _T_7155 = _T_7154 | _T_7108; // @[Mux.scala 19:72:@5511.4]
  assign _T_7156 = _T_7155 | _T_7117; // @[Mux.scala 19:72:@5512.4]
  assign _T_7157 = _T_7156 | _T_7126; // @[Mux.scala 19:72:@5513.4]
  assign _T_7158 = _T_7157 | _T_7135; // @[Mux.scala 19:72:@5514.4]
  assign _T_7159 = _T_7158 | _T_7144; // @[Mux.scala 19:72:@5515.4]
  assign _T_7160 = _T_7159 | _T_7153; // @[Mux.scala 19:72:@5516.4]
  assign _T_7402 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0}; // @[Mux.scala 19:72:@5634.4]
  assign _T_7404 = _T_1537 ? _T_7402 : 8'h0; // @[Mux.scala 19:72:@5635.4]
  assign _T_7411 = {conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1}; // @[Mux.scala 19:72:@5642.4]
  assign _T_7413 = _T_1538 ? _T_7411 : 8'h0; // @[Mux.scala 19:72:@5643.4]
  assign _T_7420 = {conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2}; // @[Mux.scala 19:72:@5650.4]
  assign _T_7422 = _T_1539 ? _T_7420 : 8'h0; // @[Mux.scala 19:72:@5651.4]
  assign _T_7429 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3}; // @[Mux.scala 19:72:@5658.4]
  assign _T_7431 = _T_1540 ? _T_7429 : 8'h0; // @[Mux.scala 19:72:@5659.4]
  assign _T_7438 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4}; // @[Mux.scala 19:72:@5666.4]
  assign _T_7440 = _T_1541 ? _T_7438 : 8'h0; // @[Mux.scala 19:72:@5667.4]
  assign _T_7447 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5}; // @[Mux.scala 19:72:@5674.4]
  assign _T_7449 = _T_1542 ? _T_7447 : 8'h0; // @[Mux.scala 19:72:@5675.4]
  assign _T_7456 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6}; // @[Mux.scala 19:72:@5682.4]
  assign _T_7458 = _T_1543 ? _T_7456 : 8'h0; // @[Mux.scala 19:72:@5683.4]
  assign _T_7465 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7}; // @[Mux.scala 19:72:@5690.4]
  assign _T_7467 = _T_1544 ? _T_7465 : 8'h0; // @[Mux.scala 19:72:@5691.4]
  assign _T_7468 = _T_7404 | _T_7413; // @[Mux.scala 19:72:@5692.4]
  assign _T_7469 = _T_7468 | _T_7422; // @[Mux.scala 19:72:@5693.4]
  assign _T_7470 = _T_7469 | _T_7431; // @[Mux.scala 19:72:@5694.4]
  assign _T_7471 = _T_7470 | _T_7440; // @[Mux.scala 19:72:@5695.4]
  assign _T_7472 = _T_7471 | _T_7449; // @[Mux.scala 19:72:@5696.4]
  assign _T_7473 = _T_7472 | _T_7458; // @[Mux.scala 19:72:@5697.4]
  assign _T_7474 = _T_7473 | _T_7467; // @[Mux.scala 19:72:@5698.4]
  assign _T_7716 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0}; // @[Mux.scala 19:72:@5816.4]
  assign _T_7718 = _T_1537 ? _T_7716 : 8'h0; // @[Mux.scala 19:72:@5817.4]
  assign _T_7725 = {conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1}; // @[Mux.scala 19:72:@5824.4]
  assign _T_7727 = _T_1538 ? _T_7725 : 8'h0; // @[Mux.scala 19:72:@5825.4]
  assign _T_7734 = {conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2}; // @[Mux.scala 19:72:@5832.4]
  assign _T_7736 = _T_1539 ? _T_7734 : 8'h0; // @[Mux.scala 19:72:@5833.4]
  assign _T_7743 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3}; // @[Mux.scala 19:72:@5840.4]
  assign _T_7745 = _T_1540 ? _T_7743 : 8'h0; // @[Mux.scala 19:72:@5841.4]
  assign _T_7752 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4}; // @[Mux.scala 19:72:@5848.4]
  assign _T_7754 = _T_1541 ? _T_7752 : 8'h0; // @[Mux.scala 19:72:@5849.4]
  assign _T_7761 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5}; // @[Mux.scala 19:72:@5856.4]
  assign _T_7763 = _T_1542 ? _T_7761 : 8'h0; // @[Mux.scala 19:72:@5857.4]
  assign _T_7770 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6}; // @[Mux.scala 19:72:@5864.4]
  assign _T_7772 = _T_1543 ? _T_7770 : 8'h0; // @[Mux.scala 19:72:@5865.4]
  assign _T_7779 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7}; // @[Mux.scala 19:72:@5872.4]
  assign _T_7781 = _T_1544 ? _T_7779 : 8'h0; // @[Mux.scala 19:72:@5873.4]
  assign _T_7782 = _T_7718 | _T_7727; // @[Mux.scala 19:72:@5874.4]
  assign _T_7783 = _T_7782 | _T_7736; // @[Mux.scala 19:72:@5875.4]
  assign _T_7784 = _T_7783 | _T_7745; // @[Mux.scala 19:72:@5876.4]
  assign _T_7785 = _T_7784 | _T_7754; // @[Mux.scala 19:72:@5877.4]
  assign _T_7786 = _T_7785 | _T_7763; // @[Mux.scala 19:72:@5878.4]
  assign _T_7787 = _T_7786 | _T_7772; // @[Mux.scala 19:72:@5879.4]
  assign _T_7788 = _T_7787 | _T_7781; // @[Mux.scala 19:72:@5880.4]
  assign _T_8030 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0}; // @[Mux.scala 19:72:@5998.4]
  assign _T_8032 = _T_1537 ? _T_8030 : 8'h0; // @[Mux.scala 19:72:@5999.4]
  assign _T_8039 = {conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1}; // @[Mux.scala 19:72:@6006.4]
  assign _T_8041 = _T_1538 ? _T_8039 : 8'h0; // @[Mux.scala 19:72:@6007.4]
  assign _T_8048 = {conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2}; // @[Mux.scala 19:72:@6014.4]
  assign _T_8050 = _T_1539 ? _T_8048 : 8'h0; // @[Mux.scala 19:72:@6015.4]
  assign _T_8057 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3}; // @[Mux.scala 19:72:@6022.4]
  assign _T_8059 = _T_1540 ? _T_8057 : 8'h0; // @[Mux.scala 19:72:@6023.4]
  assign _T_8066 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4}; // @[Mux.scala 19:72:@6030.4]
  assign _T_8068 = _T_1541 ? _T_8066 : 8'h0; // @[Mux.scala 19:72:@6031.4]
  assign _T_8075 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5}; // @[Mux.scala 19:72:@6038.4]
  assign _T_8077 = _T_1542 ? _T_8075 : 8'h0; // @[Mux.scala 19:72:@6039.4]
  assign _T_8084 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6}; // @[Mux.scala 19:72:@6046.4]
  assign _T_8086 = _T_1543 ? _T_8084 : 8'h0; // @[Mux.scala 19:72:@6047.4]
  assign _T_8093 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7}; // @[Mux.scala 19:72:@6054.4]
  assign _T_8095 = _T_1544 ? _T_8093 : 8'h0; // @[Mux.scala 19:72:@6055.4]
  assign _T_8096 = _T_8032 | _T_8041; // @[Mux.scala 19:72:@6056.4]
  assign _T_8097 = _T_8096 | _T_8050; // @[Mux.scala 19:72:@6057.4]
  assign _T_8098 = _T_8097 | _T_8059; // @[Mux.scala 19:72:@6058.4]
  assign _T_8099 = _T_8098 | _T_8068; // @[Mux.scala 19:72:@6059.4]
  assign _T_8100 = _T_8099 | _T_8077; // @[Mux.scala 19:72:@6060.4]
  assign _T_8101 = _T_8100 | _T_8086; // @[Mux.scala 19:72:@6061.4]
  assign _T_8102 = _T_8101 | _T_8095; // @[Mux.scala 19:72:@6062.4]
  assign _T_8344 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0}; // @[Mux.scala 19:72:@6180.4]
  assign _T_8346 = _T_1537 ? _T_8344 : 8'h0; // @[Mux.scala 19:72:@6181.4]
  assign _T_8353 = {conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1}; // @[Mux.scala 19:72:@6188.4]
  assign _T_8355 = _T_1538 ? _T_8353 : 8'h0; // @[Mux.scala 19:72:@6189.4]
  assign _T_8362 = {conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2}; // @[Mux.scala 19:72:@6196.4]
  assign _T_8364 = _T_1539 ? _T_8362 : 8'h0; // @[Mux.scala 19:72:@6197.4]
  assign _T_8371 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3}; // @[Mux.scala 19:72:@6204.4]
  assign _T_8373 = _T_1540 ? _T_8371 : 8'h0; // @[Mux.scala 19:72:@6205.4]
  assign _T_8380 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4}; // @[Mux.scala 19:72:@6212.4]
  assign _T_8382 = _T_1541 ? _T_8380 : 8'h0; // @[Mux.scala 19:72:@6213.4]
  assign _T_8389 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5}; // @[Mux.scala 19:72:@6220.4]
  assign _T_8391 = _T_1542 ? _T_8389 : 8'h0; // @[Mux.scala 19:72:@6221.4]
  assign _T_8398 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6}; // @[Mux.scala 19:72:@6228.4]
  assign _T_8400 = _T_1543 ? _T_8398 : 8'h0; // @[Mux.scala 19:72:@6229.4]
  assign _T_8407 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7}; // @[Mux.scala 19:72:@6236.4]
  assign _T_8409 = _T_1544 ? _T_8407 : 8'h0; // @[Mux.scala 19:72:@6237.4]
  assign _T_8410 = _T_8346 | _T_8355; // @[Mux.scala 19:72:@6238.4]
  assign _T_8411 = _T_8410 | _T_8364; // @[Mux.scala 19:72:@6239.4]
  assign _T_8412 = _T_8411 | _T_8373; // @[Mux.scala 19:72:@6240.4]
  assign _T_8413 = _T_8412 | _T_8382; // @[Mux.scala 19:72:@6241.4]
  assign _T_8414 = _T_8413 | _T_8391; // @[Mux.scala 19:72:@6242.4]
  assign _T_8415 = _T_8414 | _T_8400; // @[Mux.scala 19:72:@6243.4]
  assign _T_8416 = _T_8415 | _T_8409; // @[Mux.scala 19:72:@6244.4]
  assign _T_14526 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0}; // @[Mux.scala 19:72:@6492.4]
  assign _T_14528 = _T_1537 ? _T_14526 : 8'h0; // @[Mux.scala 19:72:@6493.4]
  assign _T_14535 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1}; // @[Mux.scala 19:72:@6500.4]
  assign _T_14537 = _T_1538 ? _T_14535 : 8'h0; // @[Mux.scala 19:72:@6501.4]
  assign _T_14544 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2}; // @[Mux.scala 19:72:@6508.4]
  assign _T_14546 = _T_1539 ? _T_14544 : 8'h0; // @[Mux.scala 19:72:@6509.4]
  assign _T_14553 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3}; // @[Mux.scala 19:72:@6516.4]
  assign _T_14555 = _T_1540 ? _T_14553 : 8'h0; // @[Mux.scala 19:72:@6517.4]
  assign _T_14562 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4}; // @[Mux.scala 19:72:@6524.4]
  assign _T_14564 = _T_1541 ? _T_14562 : 8'h0; // @[Mux.scala 19:72:@6525.4]
  assign _T_14571 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5}; // @[Mux.scala 19:72:@6532.4]
  assign _T_14573 = _T_1542 ? _T_14571 : 8'h0; // @[Mux.scala 19:72:@6533.4]
  assign _T_14580 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6}; // @[Mux.scala 19:72:@6540.4]
  assign _T_14582 = _T_1543 ? _T_14580 : 8'h0; // @[Mux.scala 19:72:@6541.4]
  assign _T_14589 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7}; // @[Mux.scala 19:72:@6548.4]
  assign _T_14591 = _T_1544 ? _T_14589 : 8'h0; // @[Mux.scala 19:72:@6549.4]
  assign _T_14592 = _T_14528 | _T_14537; // @[Mux.scala 19:72:@6550.4]
  assign _T_14593 = _T_14592 | _T_14546; // @[Mux.scala 19:72:@6551.4]
  assign _T_14594 = _T_14593 | _T_14555; // @[Mux.scala 19:72:@6552.4]
  assign _T_14595 = _T_14594 | _T_14564; // @[Mux.scala 19:72:@6553.4]
  assign _T_14596 = _T_14595 | _T_14573; // @[Mux.scala 19:72:@6554.4]
  assign _T_14597 = _T_14596 | _T_14582; // @[Mux.scala 19:72:@6555.4]
  assign _T_14598 = _T_14597 | _T_14591; // @[Mux.scala 19:72:@6556.4]
  assign _T_14840 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0}; // @[Mux.scala 19:72:@6674.4]
  assign _T_14842 = _T_1537 ? _T_14840 : 8'h0; // @[Mux.scala 19:72:@6675.4]
  assign _T_14849 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1}; // @[Mux.scala 19:72:@6682.4]
  assign _T_14851 = _T_1538 ? _T_14849 : 8'h0; // @[Mux.scala 19:72:@6683.4]
  assign _T_14858 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2}; // @[Mux.scala 19:72:@6690.4]
  assign _T_14860 = _T_1539 ? _T_14858 : 8'h0; // @[Mux.scala 19:72:@6691.4]
  assign _T_14867 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3}; // @[Mux.scala 19:72:@6698.4]
  assign _T_14869 = _T_1540 ? _T_14867 : 8'h0; // @[Mux.scala 19:72:@6699.4]
  assign _T_14876 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4}; // @[Mux.scala 19:72:@6706.4]
  assign _T_14878 = _T_1541 ? _T_14876 : 8'h0; // @[Mux.scala 19:72:@6707.4]
  assign _T_14885 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5}; // @[Mux.scala 19:72:@6714.4]
  assign _T_14887 = _T_1542 ? _T_14885 : 8'h0; // @[Mux.scala 19:72:@6715.4]
  assign _T_14894 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6}; // @[Mux.scala 19:72:@6722.4]
  assign _T_14896 = _T_1543 ? _T_14894 : 8'h0; // @[Mux.scala 19:72:@6723.4]
  assign _T_14903 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7}; // @[Mux.scala 19:72:@6730.4]
  assign _T_14905 = _T_1544 ? _T_14903 : 8'h0; // @[Mux.scala 19:72:@6731.4]
  assign _T_14906 = _T_14842 | _T_14851; // @[Mux.scala 19:72:@6732.4]
  assign _T_14907 = _T_14906 | _T_14860; // @[Mux.scala 19:72:@6733.4]
  assign _T_14908 = _T_14907 | _T_14869; // @[Mux.scala 19:72:@6734.4]
  assign _T_14909 = _T_14908 | _T_14878; // @[Mux.scala 19:72:@6735.4]
  assign _T_14910 = _T_14909 | _T_14887; // @[Mux.scala 19:72:@6736.4]
  assign _T_14911 = _T_14910 | _T_14896; // @[Mux.scala 19:72:@6737.4]
  assign _T_14912 = _T_14911 | _T_14905; // @[Mux.scala 19:72:@6738.4]
  assign _T_15154 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0}; // @[Mux.scala 19:72:@6856.4]
  assign _T_15156 = _T_1537 ? _T_15154 : 8'h0; // @[Mux.scala 19:72:@6857.4]
  assign _T_15163 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1}; // @[Mux.scala 19:72:@6864.4]
  assign _T_15165 = _T_1538 ? _T_15163 : 8'h0; // @[Mux.scala 19:72:@6865.4]
  assign _T_15172 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2}; // @[Mux.scala 19:72:@6872.4]
  assign _T_15174 = _T_1539 ? _T_15172 : 8'h0; // @[Mux.scala 19:72:@6873.4]
  assign _T_15181 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3}; // @[Mux.scala 19:72:@6880.4]
  assign _T_15183 = _T_1540 ? _T_15181 : 8'h0; // @[Mux.scala 19:72:@6881.4]
  assign _T_15190 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4}; // @[Mux.scala 19:72:@6888.4]
  assign _T_15192 = _T_1541 ? _T_15190 : 8'h0; // @[Mux.scala 19:72:@6889.4]
  assign _T_15199 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5}; // @[Mux.scala 19:72:@6896.4]
  assign _T_15201 = _T_1542 ? _T_15199 : 8'h0; // @[Mux.scala 19:72:@6897.4]
  assign _T_15208 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6}; // @[Mux.scala 19:72:@6904.4]
  assign _T_15210 = _T_1543 ? _T_15208 : 8'h0; // @[Mux.scala 19:72:@6905.4]
  assign _T_15217 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7}; // @[Mux.scala 19:72:@6912.4]
  assign _T_15219 = _T_1544 ? _T_15217 : 8'h0; // @[Mux.scala 19:72:@6913.4]
  assign _T_15220 = _T_15156 | _T_15165; // @[Mux.scala 19:72:@6914.4]
  assign _T_15221 = _T_15220 | _T_15174; // @[Mux.scala 19:72:@6915.4]
  assign _T_15222 = _T_15221 | _T_15183; // @[Mux.scala 19:72:@6916.4]
  assign _T_15223 = _T_15222 | _T_15192; // @[Mux.scala 19:72:@6917.4]
  assign _T_15224 = _T_15223 | _T_15201; // @[Mux.scala 19:72:@6918.4]
  assign _T_15225 = _T_15224 | _T_15210; // @[Mux.scala 19:72:@6919.4]
  assign _T_15226 = _T_15225 | _T_15219; // @[Mux.scala 19:72:@6920.4]
  assign _T_15468 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0}; // @[Mux.scala 19:72:@7038.4]
  assign _T_15470 = _T_1537 ? _T_15468 : 8'h0; // @[Mux.scala 19:72:@7039.4]
  assign _T_15477 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1}; // @[Mux.scala 19:72:@7046.4]
  assign _T_15479 = _T_1538 ? _T_15477 : 8'h0; // @[Mux.scala 19:72:@7047.4]
  assign _T_15486 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2}; // @[Mux.scala 19:72:@7054.4]
  assign _T_15488 = _T_1539 ? _T_15486 : 8'h0; // @[Mux.scala 19:72:@7055.4]
  assign _T_15495 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3}; // @[Mux.scala 19:72:@7062.4]
  assign _T_15497 = _T_1540 ? _T_15495 : 8'h0; // @[Mux.scala 19:72:@7063.4]
  assign _T_15504 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4}; // @[Mux.scala 19:72:@7070.4]
  assign _T_15506 = _T_1541 ? _T_15504 : 8'h0; // @[Mux.scala 19:72:@7071.4]
  assign _T_15513 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5}; // @[Mux.scala 19:72:@7078.4]
  assign _T_15515 = _T_1542 ? _T_15513 : 8'h0; // @[Mux.scala 19:72:@7079.4]
  assign _T_15522 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6}; // @[Mux.scala 19:72:@7086.4]
  assign _T_15524 = _T_1543 ? _T_15522 : 8'h0; // @[Mux.scala 19:72:@7087.4]
  assign _T_15531 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7}; // @[Mux.scala 19:72:@7094.4]
  assign _T_15533 = _T_1544 ? _T_15531 : 8'h0; // @[Mux.scala 19:72:@7095.4]
  assign _T_15534 = _T_15470 | _T_15479; // @[Mux.scala 19:72:@7096.4]
  assign _T_15535 = _T_15534 | _T_15488; // @[Mux.scala 19:72:@7097.4]
  assign _T_15536 = _T_15535 | _T_15497; // @[Mux.scala 19:72:@7098.4]
  assign _T_15537 = _T_15536 | _T_15506; // @[Mux.scala 19:72:@7099.4]
  assign _T_15538 = _T_15537 | _T_15515; // @[Mux.scala 19:72:@7100.4]
  assign _T_15539 = _T_15538 | _T_15524; // @[Mux.scala 19:72:@7101.4]
  assign _T_15540 = _T_15539 | _T_15533; // @[Mux.scala 19:72:@7102.4]
  assign _T_15782 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0}; // @[Mux.scala 19:72:@7220.4]
  assign _T_15784 = _T_1537 ? _T_15782 : 8'h0; // @[Mux.scala 19:72:@7221.4]
  assign _T_15791 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1}; // @[Mux.scala 19:72:@7228.4]
  assign _T_15793 = _T_1538 ? _T_15791 : 8'h0; // @[Mux.scala 19:72:@7229.4]
  assign _T_15800 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2}; // @[Mux.scala 19:72:@7236.4]
  assign _T_15802 = _T_1539 ? _T_15800 : 8'h0; // @[Mux.scala 19:72:@7237.4]
  assign _T_15809 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3}; // @[Mux.scala 19:72:@7244.4]
  assign _T_15811 = _T_1540 ? _T_15809 : 8'h0; // @[Mux.scala 19:72:@7245.4]
  assign _T_15818 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4}; // @[Mux.scala 19:72:@7252.4]
  assign _T_15820 = _T_1541 ? _T_15818 : 8'h0; // @[Mux.scala 19:72:@7253.4]
  assign _T_15827 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5}; // @[Mux.scala 19:72:@7260.4]
  assign _T_15829 = _T_1542 ? _T_15827 : 8'h0; // @[Mux.scala 19:72:@7261.4]
  assign _T_15836 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6}; // @[Mux.scala 19:72:@7268.4]
  assign _T_15838 = _T_1543 ? _T_15836 : 8'h0; // @[Mux.scala 19:72:@7269.4]
  assign _T_15845 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7}; // @[Mux.scala 19:72:@7276.4]
  assign _T_15847 = _T_1544 ? _T_15845 : 8'h0; // @[Mux.scala 19:72:@7277.4]
  assign _T_15848 = _T_15784 | _T_15793; // @[Mux.scala 19:72:@7278.4]
  assign _T_15849 = _T_15848 | _T_15802; // @[Mux.scala 19:72:@7279.4]
  assign _T_15850 = _T_15849 | _T_15811; // @[Mux.scala 19:72:@7280.4]
  assign _T_15851 = _T_15850 | _T_15820; // @[Mux.scala 19:72:@7281.4]
  assign _T_15852 = _T_15851 | _T_15829; // @[Mux.scala 19:72:@7282.4]
  assign _T_15853 = _T_15852 | _T_15838; // @[Mux.scala 19:72:@7283.4]
  assign _T_15854 = _T_15853 | _T_15847; // @[Mux.scala 19:72:@7284.4]
  assign _T_16096 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0}; // @[Mux.scala 19:72:@7402.4]
  assign _T_16098 = _T_1537 ? _T_16096 : 8'h0; // @[Mux.scala 19:72:@7403.4]
  assign _T_16105 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1}; // @[Mux.scala 19:72:@7410.4]
  assign _T_16107 = _T_1538 ? _T_16105 : 8'h0; // @[Mux.scala 19:72:@7411.4]
  assign _T_16114 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2}; // @[Mux.scala 19:72:@7418.4]
  assign _T_16116 = _T_1539 ? _T_16114 : 8'h0; // @[Mux.scala 19:72:@7419.4]
  assign _T_16123 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3}; // @[Mux.scala 19:72:@7426.4]
  assign _T_16125 = _T_1540 ? _T_16123 : 8'h0; // @[Mux.scala 19:72:@7427.4]
  assign _T_16132 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4}; // @[Mux.scala 19:72:@7434.4]
  assign _T_16134 = _T_1541 ? _T_16132 : 8'h0; // @[Mux.scala 19:72:@7435.4]
  assign _T_16141 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5}; // @[Mux.scala 19:72:@7442.4]
  assign _T_16143 = _T_1542 ? _T_16141 : 8'h0; // @[Mux.scala 19:72:@7443.4]
  assign _T_16150 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6}; // @[Mux.scala 19:72:@7450.4]
  assign _T_16152 = _T_1543 ? _T_16150 : 8'h0; // @[Mux.scala 19:72:@7451.4]
  assign _T_16159 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7}; // @[Mux.scala 19:72:@7458.4]
  assign _T_16161 = _T_1544 ? _T_16159 : 8'h0; // @[Mux.scala 19:72:@7459.4]
  assign _T_16162 = _T_16098 | _T_16107; // @[Mux.scala 19:72:@7460.4]
  assign _T_16163 = _T_16162 | _T_16116; // @[Mux.scala 19:72:@7461.4]
  assign _T_16164 = _T_16163 | _T_16125; // @[Mux.scala 19:72:@7462.4]
  assign _T_16165 = _T_16164 | _T_16134; // @[Mux.scala 19:72:@7463.4]
  assign _T_16166 = _T_16165 | _T_16143; // @[Mux.scala 19:72:@7464.4]
  assign _T_16167 = _T_16166 | _T_16152; // @[Mux.scala 19:72:@7465.4]
  assign _T_16168 = _T_16167 | _T_16161; // @[Mux.scala 19:72:@7466.4]
  assign _T_16410 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0}; // @[Mux.scala 19:72:@7584.4]
  assign _T_16412 = _T_1537 ? _T_16410 : 8'h0; // @[Mux.scala 19:72:@7585.4]
  assign _T_16419 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1}; // @[Mux.scala 19:72:@7592.4]
  assign _T_16421 = _T_1538 ? _T_16419 : 8'h0; // @[Mux.scala 19:72:@7593.4]
  assign _T_16428 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2}; // @[Mux.scala 19:72:@7600.4]
  assign _T_16430 = _T_1539 ? _T_16428 : 8'h0; // @[Mux.scala 19:72:@7601.4]
  assign _T_16437 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3}; // @[Mux.scala 19:72:@7608.4]
  assign _T_16439 = _T_1540 ? _T_16437 : 8'h0; // @[Mux.scala 19:72:@7609.4]
  assign _T_16446 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4}; // @[Mux.scala 19:72:@7616.4]
  assign _T_16448 = _T_1541 ? _T_16446 : 8'h0; // @[Mux.scala 19:72:@7617.4]
  assign _T_16455 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5}; // @[Mux.scala 19:72:@7624.4]
  assign _T_16457 = _T_1542 ? _T_16455 : 8'h0; // @[Mux.scala 19:72:@7625.4]
  assign _T_16464 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6}; // @[Mux.scala 19:72:@7632.4]
  assign _T_16466 = _T_1543 ? _T_16464 : 8'h0; // @[Mux.scala 19:72:@7633.4]
  assign _T_16473 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7}; // @[Mux.scala 19:72:@7640.4]
  assign _T_16475 = _T_1544 ? _T_16473 : 8'h0; // @[Mux.scala 19:72:@7641.4]
  assign _T_16476 = _T_16412 | _T_16421; // @[Mux.scala 19:72:@7642.4]
  assign _T_16477 = _T_16476 | _T_16430; // @[Mux.scala 19:72:@7643.4]
  assign _T_16478 = _T_16477 | _T_16439; // @[Mux.scala 19:72:@7644.4]
  assign _T_16479 = _T_16478 | _T_16448; // @[Mux.scala 19:72:@7645.4]
  assign _T_16480 = _T_16479 | _T_16457; // @[Mux.scala 19:72:@7646.4]
  assign _T_16481 = _T_16480 | _T_16466; // @[Mux.scala 19:72:@7647.4]
  assign _T_16482 = _T_16481 | _T_16475; // @[Mux.scala 19:72:@7648.4]
  assign _T_16724 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0}; // @[Mux.scala 19:72:@7766.4]
  assign _T_16726 = _T_1537 ? _T_16724 : 8'h0; // @[Mux.scala 19:72:@7767.4]
  assign _T_16733 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1}; // @[Mux.scala 19:72:@7774.4]
  assign _T_16735 = _T_1538 ? _T_16733 : 8'h0; // @[Mux.scala 19:72:@7775.4]
  assign _T_16742 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2}; // @[Mux.scala 19:72:@7782.4]
  assign _T_16744 = _T_1539 ? _T_16742 : 8'h0; // @[Mux.scala 19:72:@7783.4]
  assign _T_16751 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3}; // @[Mux.scala 19:72:@7790.4]
  assign _T_16753 = _T_1540 ? _T_16751 : 8'h0; // @[Mux.scala 19:72:@7791.4]
  assign _T_16760 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4}; // @[Mux.scala 19:72:@7798.4]
  assign _T_16762 = _T_1541 ? _T_16760 : 8'h0; // @[Mux.scala 19:72:@7799.4]
  assign _T_16769 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5}; // @[Mux.scala 19:72:@7806.4]
  assign _T_16771 = _T_1542 ? _T_16769 : 8'h0; // @[Mux.scala 19:72:@7807.4]
  assign _T_16778 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6}; // @[Mux.scala 19:72:@7814.4]
  assign _T_16780 = _T_1543 ? _T_16778 : 8'h0; // @[Mux.scala 19:72:@7815.4]
  assign _T_16787 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7}; // @[Mux.scala 19:72:@7822.4]
  assign _T_16789 = _T_1544 ? _T_16787 : 8'h0; // @[Mux.scala 19:72:@7823.4]
  assign _T_16790 = _T_16726 | _T_16735; // @[Mux.scala 19:72:@7824.4]
  assign _T_16791 = _T_16790 | _T_16744; // @[Mux.scala 19:72:@7825.4]
  assign _T_16792 = _T_16791 | _T_16753; // @[Mux.scala 19:72:@7826.4]
  assign _T_16793 = _T_16792 | _T_16762; // @[Mux.scala 19:72:@7827.4]
  assign _T_16794 = _T_16793 | _T_16771; // @[Mux.scala 19:72:@7828.4]
  assign _T_16795 = _T_16794 | _T_16780; // @[Mux.scala 19:72:@7829.4]
  assign _T_16796 = _T_16795 | _T_16789; // @[Mux.scala 19:72:@7830.4]
  assign _T_23556 = conflictPReg_0_2 ? 2'h2 : {{1'd0}, conflictPReg_0_1}; // @[LoadQueue.scala 191:60:@8047.4]
  assign _T_23557 = conflictPReg_0_3 ? 2'h3 : _T_23556; // @[LoadQueue.scala 191:60:@8048.4]
  assign _T_23558 = conflictPReg_0_4 ? 3'h4 : {{1'd0}, _T_23557}; // @[LoadQueue.scala 191:60:@8049.4]
  assign _T_23559 = conflictPReg_0_5 ? 3'h5 : _T_23558; // @[LoadQueue.scala 191:60:@8050.4]
  assign _T_23560 = conflictPReg_0_6 ? 3'h6 : _T_23559; // @[LoadQueue.scala 191:60:@8051.4]
  assign _T_23561 = conflictPReg_0_7 ? 3'h7 : _T_23560; // @[LoadQueue.scala 191:60:@8052.4]
  assign _T_23564 = conflictPReg_0_0 | conflictPReg_0_1; // @[LoadQueue.scala 192:43:@8054.4]
  assign _T_23565 = _T_23564 | conflictPReg_0_2; // @[LoadQueue.scala 192:43:@8055.4]
  assign _T_23566 = _T_23565 | conflictPReg_0_3; // @[LoadQueue.scala 192:43:@8056.4]
  assign _T_23567 = _T_23566 | conflictPReg_0_4; // @[LoadQueue.scala 192:43:@8057.4]
  assign _T_23568 = _T_23567 | conflictPReg_0_5; // @[LoadQueue.scala 192:43:@8058.4]
  assign _T_23569 = _T_23568 | conflictPReg_0_6; // @[LoadQueue.scala 192:43:@8059.4]
  assign _T_23570 = _T_23569 | conflictPReg_0_7; // @[LoadQueue.scala 192:43:@8060.4]
  assign _GEN_240 = 3'h0 == _T_23561; // @[LoadQueue.scala 193:43:@8062.6]
  assign _GEN_241 = 3'h1 == _T_23561; // @[LoadQueue.scala 193:43:@8062.6]
  assign _GEN_242 = 3'h2 == _T_23561; // @[LoadQueue.scala 193:43:@8062.6]
  assign _GEN_243 = 3'h3 == _T_23561; // @[LoadQueue.scala 193:43:@8062.6]
  assign _GEN_244 = 3'h4 == _T_23561; // @[LoadQueue.scala 193:43:@8062.6]
  assign _GEN_245 = 3'h5 == _T_23561; // @[LoadQueue.scala 193:43:@8062.6]
  assign _GEN_246 = 3'h6 == _T_23561; // @[LoadQueue.scala 193:43:@8062.6]
  assign _GEN_247 = 3'h7 == _T_23561; // @[LoadQueue.scala 193:43:@8062.6]
  assign _GEN_249 = 3'h1 == _T_23561 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8063.6]
  assign _GEN_250 = 3'h2 == _T_23561 ? shiftedStoreDataKnownPReg_2 : _GEN_249; // @[LoadQueue.scala 194:31:@8063.6]
  assign _GEN_251 = 3'h3 == _T_23561 ? shiftedStoreDataKnownPReg_3 : _GEN_250; // @[LoadQueue.scala 194:31:@8063.6]
  assign _GEN_252 = 3'h4 == _T_23561 ? shiftedStoreDataKnownPReg_4 : _GEN_251; // @[LoadQueue.scala 194:31:@8063.6]
  assign _GEN_253 = 3'h5 == _T_23561 ? shiftedStoreDataKnownPReg_5 : _GEN_252; // @[LoadQueue.scala 194:31:@8063.6]
  assign _GEN_254 = 3'h6 == _T_23561 ? shiftedStoreDataKnownPReg_6 : _GEN_253; // @[LoadQueue.scala 194:31:@8063.6]
  assign _GEN_255 = 3'h7 == _T_23561 ? shiftedStoreDataKnownPReg_7 : _GEN_254; // @[LoadQueue.scala 194:31:@8063.6]
  assign _GEN_257 = 3'h1 == _T_23561 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8064.6]
  assign _GEN_258 = 3'h2 == _T_23561 ? shiftedStoreDataQPreg_2 : _GEN_257; // @[LoadQueue.scala 195:31:@8064.6]
  assign _GEN_259 = 3'h3 == _T_23561 ? shiftedStoreDataQPreg_3 : _GEN_258; // @[LoadQueue.scala 195:31:@8064.6]
  assign _GEN_260 = 3'h4 == _T_23561 ? shiftedStoreDataQPreg_4 : _GEN_259; // @[LoadQueue.scala 195:31:@8064.6]
  assign _GEN_261 = 3'h5 == _T_23561 ? shiftedStoreDataQPreg_5 : _GEN_260; // @[LoadQueue.scala 195:31:@8064.6]
  assign _GEN_262 = 3'h6 == _T_23561 ? shiftedStoreDataQPreg_6 : _GEN_261; // @[LoadQueue.scala 195:31:@8064.6]
  assign _GEN_263 = 3'h7 == _T_23561 ? shiftedStoreDataQPreg_7 : _GEN_262; // @[LoadQueue.scala 195:31:@8064.6]
  assign lastConflict_0_0 = _T_23570 ? _GEN_240 : 1'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign lastConflict_0_1 = _T_23570 ? _GEN_241 : 1'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign lastConflict_0_2 = _T_23570 ? _GEN_242 : 1'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign lastConflict_0_3 = _T_23570 ? _GEN_243 : 1'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign lastConflict_0_4 = _T_23570 ? _GEN_244 : 1'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign lastConflict_0_5 = _T_23570 ? _GEN_245 : 1'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign lastConflict_0_6 = _T_23570 ? _GEN_246 : 1'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign lastConflict_0_7 = _T_23570 ? _GEN_247 : 1'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign canBypass_0 = _T_23570 ? _GEN_255 : 1'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign bypassVal_0 = _T_23570 ? _GEN_263 : 32'h0; // @[LoadQueue.scala 192:53:@8061.4]
  assign _T_23636 = conflictPReg_1_2 ? 2'h2 : {{1'd0}, conflictPReg_1_1}; // @[LoadQueue.scala 191:60:@8094.4]
  assign _T_23637 = conflictPReg_1_3 ? 2'h3 : _T_23636; // @[LoadQueue.scala 191:60:@8095.4]
  assign _T_23638 = conflictPReg_1_4 ? 3'h4 : {{1'd0}, _T_23637}; // @[LoadQueue.scala 191:60:@8096.4]
  assign _T_23639 = conflictPReg_1_5 ? 3'h5 : _T_23638; // @[LoadQueue.scala 191:60:@8097.4]
  assign _T_23640 = conflictPReg_1_6 ? 3'h6 : _T_23639; // @[LoadQueue.scala 191:60:@8098.4]
  assign _T_23641 = conflictPReg_1_7 ? 3'h7 : _T_23640; // @[LoadQueue.scala 191:60:@8099.4]
  assign _T_23644 = conflictPReg_1_0 | conflictPReg_1_1; // @[LoadQueue.scala 192:43:@8101.4]
  assign _T_23645 = _T_23644 | conflictPReg_1_2; // @[LoadQueue.scala 192:43:@8102.4]
  assign _T_23646 = _T_23645 | conflictPReg_1_3; // @[LoadQueue.scala 192:43:@8103.4]
  assign _T_23647 = _T_23646 | conflictPReg_1_4; // @[LoadQueue.scala 192:43:@8104.4]
  assign _T_23648 = _T_23647 | conflictPReg_1_5; // @[LoadQueue.scala 192:43:@8105.4]
  assign _T_23649 = _T_23648 | conflictPReg_1_6; // @[LoadQueue.scala 192:43:@8106.4]
  assign _T_23650 = _T_23649 | conflictPReg_1_7; // @[LoadQueue.scala 192:43:@8107.4]
  assign _GEN_274 = 3'h0 == _T_23641; // @[LoadQueue.scala 193:43:@8109.6]
  assign _GEN_275 = 3'h1 == _T_23641; // @[LoadQueue.scala 193:43:@8109.6]
  assign _GEN_276 = 3'h2 == _T_23641; // @[LoadQueue.scala 193:43:@8109.6]
  assign _GEN_277 = 3'h3 == _T_23641; // @[LoadQueue.scala 193:43:@8109.6]
  assign _GEN_278 = 3'h4 == _T_23641; // @[LoadQueue.scala 193:43:@8109.6]
  assign _GEN_279 = 3'h5 == _T_23641; // @[LoadQueue.scala 193:43:@8109.6]
  assign _GEN_280 = 3'h6 == _T_23641; // @[LoadQueue.scala 193:43:@8109.6]
  assign _GEN_281 = 3'h7 == _T_23641; // @[LoadQueue.scala 193:43:@8109.6]
  assign _GEN_283 = 3'h1 == _T_23641 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8110.6]
  assign _GEN_284 = 3'h2 == _T_23641 ? shiftedStoreDataKnownPReg_2 : _GEN_283; // @[LoadQueue.scala 194:31:@8110.6]
  assign _GEN_285 = 3'h3 == _T_23641 ? shiftedStoreDataKnownPReg_3 : _GEN_284; // @[LoadQueue.scala 194:31:@8110.6]
  assign _GEN_286 = 3'h4 == _T_23641 ? shiftedStoreDataKnownPReg_4 : _GEN_285; // @[LoadQueue.scala 194:31:@8110.6]
  assign _GEN_287 = 3'h5 == _T_23641 ? shiftedStoreDataKnownPReg_5 : _GEN_286; // @[LoadQueue.scala 194:31:@8110.6]
  assign _GEN_288 = 3'h6 == _T_23641 ? shiftedStoreDataKnownPReg_6 : _GEN_287; // @[LoadQueue.scala 194:31:@8110.6]
  assign _GEN_289 = 3'h7 == _T_23641 ? shiftedStoreDataKnownPReg_7 : _GEN_288; // @[LoadQueue.scala 194:31:@8110.6]
  assign _GEN_291 = 3'h1 == _T_23641 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8111.6]
  assign _GEN_292 = 3'h2 == _T_23641 ? shiftedStoreDataQPreg_2 : _GEN_291; // @[LoadQueue.scala 195:31:@8111.6]
  assign _GEN_293 = 3'h3 == _T_23641 ? shiftedStoreDataQPreg_3 : _GEN_292; // @[LoadQueue.scala 195:31:@8111.6]
  assign _GEN_294 = 3'h4 == _T_23641 ? shiftedStoreDataQPreg_4 : _GEN_293; // @[LoadQueue.scala 195:31:@8111.6]
  assign _GEN_295 = 3'h5 == _T_23641 ? shiftedStoreDataQPreg_5 : _GEN_294; // @[LoadQueue.scala 195:31:@8111.6]
  assign _GEN_296 = 3'h6 == _T_23641 ? shiftedStoreDataQPreg_6 : _GEN_295; // @[LoadQueue.scala 195:31:@8111.6]
  assign _GEN_297 = 3'h7 == _T_23641 ? shiftedStoreDataQPreg_7 : _GEN_296; // @[LoadQueue.scala 195:31:@8111.6]
  assign lastConflict_1_0 = _T_23650 ? _GEN_274 : 1'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign lastConflict_1_1 = _T_23650 ? _GEN_275 : 1'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign lastConflict_1_2 = _T_23650 ? _GEN_276 : 1'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign lastConflict_1_3 = _T_23650 ? _GEN_277 : 1'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign lastConflict_1_4 = _T_23650 ? _GEN_278 : 1'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign lastConflict_1_5 = _T_23650 ? _GEN_279 : 1'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign lastConflict_1_6 = _T_23650 ? _GEN_280 : 1'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign lastConflict_1_7 = _T_23650 ? _GEN_281 : 1'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign canBypass_1 = _T_23650 ? _GEN_289 : 1'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign bypassVal_1 = _T_23650 ? _GEN_297 : 32'h0; // @[LoadQueue.scala 192:53:@8108.4]
  assign _T_23716 = conflictPReg_2_2 ? 2'h2 : {{1'd0}, conflictPReg_2_1}; // @[LoadQueue.scala 191:60:@8141.4]
  assign _T_23717 = conflictPReg_2_3 ? 2'h3 : _T_23716; // @[LoadQueue.scala 191:60:@8142.4]
  assign _T_23718 = conflictPReg_2_4 ? 3'h4 : {{1'd0}, _T_23717}; // @[LoadQueue.scala 191:60:@8143.4]
  assign _T_23719 = conflictPReg_2_5 ? 3'h5 : _T_23718; // @[LoadQueue.scala 191:60:@8144.4]
  assign _T_23720 = conflictPReg_2_6 ? 3'h6 : _T_23719; // @[LoadQueue.scala 191:60:@8145.4]
  assign _T_23721 = conflictPReg_2_7 ? 3'h7 : _T_23720; // @[LoadQueue.scala 191:60:@8146.4]
  assign _T_23724 = conflictPReg_2_0 | conflictPReg_2_1; // @[LoadQueue.scala 192:43:@8148.4]
  assign _T_23725 = _T_23724 | conflictPReg_2_2; // @[LoadQueue.scala 192:43:@8149.4]
  assign _T_23726 = _T_23725 | conflictPReg_2_3; // @[LoadQueue.scala 192:43:@8150.4]
  assign _T_23727 = _T_23726 | conflictPReg_2_4; // @[LoadQueue.scala 192:43:@8151.4]
  assign _T_23728 = _T_23727 | conflictPReg_2_5; // @[LoadQueue.scala 192:43:@8152.4]
  assign _T_23729 = _T_23728 | conflictPReg_2_6; // @[LoadQueue.scala 192:43:@8153.4]
  assign _T_23730 = _T_23729 | conflictPReg_2_7; // @[LoadQueue.scala 192:43:@8154.4]
  assign _GEN_308 = 3'h0 == _T_23721; // @[LoadQueue.scala 193:43:@8156.6]
  assign _GEN_309 = 3'h1 == _T_23721; // @[LoadQueue.scala 193:43:@8156.6]
  assign _GEN_310 = 3'h2 == _T_23721; // @[LoadQueue.scala 193:43:@8156.6]
  assign _GEN_311 = 3'h3 == _T_23721; // @[LoadQueue.scala 193:43:@8156.6]
  assign _GEN_312 = 3'h4 == _T_23721; // @[LoadQueue.scala 193:43:@8156.6]
  assign _GEN_313 = 3'h5 == _T_23721; // @[LoadQueue.scala 193:43:@8156.6]
  assign _GEN_314 = 3'h6 == _T_23721; // @[LoadQueue.scala 193:43:@8156.6]
  assign _GEN_315 = 3'h7 == _T_23721; // @[LoadQueue.scala 193:43:@8156.6]
  assign _GEN_317 = 3'h1 == _T_23721 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8157.6]
  assign _GEN_318 = 3'h2 == _T_23721 ? shiftedStoreDataKnownPReg_2 : _GEN_317; // @[LoadQueue.scala 194:31:@8157.6]
  assign _GEN_319 = 3'h3 == _T_23721 ? shiftedStoreDataKnownPReg_3 : _GEN_318; // @[LoadQueue.scala 194:31:@8157.6]
  assign _GEN_320 = 3'h4 == _T_23721 ? shiftedStoreDataKnownPReg_4 : _GEN_319; // @[LoadQueue.scala 194:31:@8157.6]
  assign _GEN_321 = 3'h5 == _T_23721 ? shiftedStoreDataKnownPReg_5 : _GEN_320; // @[LoadQueue.scala 194:31:@8157.6]
  assign _GEN_322 = 3'h6 == _T_23721 ? shiftedStoreDataKnownPReg_6 : _GEN_321; // @[LoadQueue.scala 194:31:@8157.6]
  assign _GEN_323 = 3'h7 == _T_23721 ? shiftedStoreDataKnownPReg_7 : _GEN_322; // @[LoadQueue.scala 194:31:@8157.6]
  assign _GEN_325 = 3'h1 == _T_23721 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8158.6]
  assign _GEN_326 = 3'h2 == _T_23721 ? shiftedStoreDataQPreg_2 : _GEN_325; // @[LoadQueue.scala 195:31:@8158.6]
  assign _GEN_327 = 3'h3 == _T_23721 ? shiftedStoreDataQPreg_3 : _GEN_326; // @[LoadQueue.scala 195:31:@8158.6]
  assign _GEN_328 = 3'h4 == _T_23721 ? shiftedStoreDataQPreg_4 : _GEN_327; // @[LoadQueue.scala 195:31:@8158.6]
  assign _GEN_329 = 3'h5 == _T_23721 ? shiftedStoreDataQPreg_5 : _GEN_328; // @[LoadQueue.scala 195:31:@8158.6]
  assign _GEN_330 = 3'h6 == _T_23721 ? shiftedStoreDataQPreg_6 : _GEN_329; // @[LoadQueue.scala 195:31:@8158.6]
  assign _GEN_331 = 3'h7 == _T_23721 ? shiftedStoreDataQPreg_7 : _GEN_330; // @[LoadQueue.scala 195:31:@8158.6]
  assign lastConflict_2_0 = _T_23730 ? _GEN_308 : 1'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign lastConflict_2_1 = _T_23730 ? _GEN_309 : 1'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign lastConflict_2_2 = _T_23730 ? _GEN_310 : 1'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign lastConflict_2_3 = _T_23730 ? _GEN_311 : 1'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign lastConflict_2_4 = _T_23730 ? _GEN_312 : 1'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign lastConflict_2_5 = _T_23730 ? _GEN_313 : 1'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign lastConflict_2_6 = _T_23730 ? _GEN_314 : 1'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign lastConflict_2_7 = _T_23730 ? _GEN_315 : 1'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign canBypass_2 = _T_23730 ? _GEN_323 : 1'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign bypassVal_2 = _T_23730 ? _GEN_331 : 32'h0; // @[LoadQueue.scala 192:53:@8155.4]
  assign _T_23796 = conflictPReg_3_2 ? 2'h2 : {{1'd0}, conflictPReg_3_1}; // @[LoadQueue.scala 191:60:@8188.4]
  assign _T_23797 = conflictPReg_3_3 ? 2'h3 : _T_23796; // @[LoadQueue.scala 191:60:@8189.4]
  assign _T_23798 = conflictPReg_3_4 ? 3'h4 : {{1'd0}, _T_23797}; // @[LoadQueue.scala 191:60:@8190.4]
  assign _T_23799 = conflictPReg_3_5 ? 3'h5 : _T_23798; // @[LoadQueue.scala 191:60:@8191.4]
  assign _T_23800 = conflictPReg_3_6 ? 3'h6 : _T_23799; // @[LoadQueue.scala 191:60:@8192.4]
  assign _T_23801 = conflictPReg_3_7 ? 3'h7 : _T_23800; // @[LoadQueue.scala 191:60:@8193.4]
  assign _T_23804 = conflictPReg_3_0 | conflictPReg_3_1; // @[LoadQueue.scala 192:43:@8195.4]
  assign _T_23805 = _T_23804 | conflictPReg_3_2; // @[LoadQueue.scala 192:43:@8196.4]
  assign _T_23806 = _T_23805 | conflictPReg_3_3; // @[LoadQueue.scala 192:43:@8197.4]
  assign _T_23807 = _T_23806 | conflictPReg_3_4; // @[LoadQueue.scala 192:43:@8198.4]
  assign _T_23808 = _T_23807 | conflictPReg_3_5; // @[LoadQueue.scala 192:43:@8199.4]
  assign _T_23809 = _T_23808 | conflictPReg_3_6; // @[LoadQueue.scala 192:43:@8200.4]
  assign _T_23810 = _T_23809 | conflictPReg_3_7; // @[LoadQueue.scala 192:43:@8201.4]
  assign _GEN_342 = 3'h0 == _T_23801; // @[LoadQueue.scala 193:43:@8203.6]
  assign _GEN_343 = 3'h1 == _T_23801; // @[LoadQueue.scala 193:43:@8203.6]
  assign _GEN_344 = 3'h2 == _T_23801; // @[LoadQueue.scala 193:43:@8203.6]
  assign _GEN_345 = 3'h3 == _T_23801; // @[LoadQueue.scala 193:43:@8203.6]
  assign _GEN_346 = 3'h4 == _T_23801; // @[LoadQueue.scala 193:43:@8203.6]
  assign _GEN_347 = 3'h5 == _T_23801; // @[LoadQueue.scala 193:43:@8203.6]
  assign _GEN_348 = 3'h6 == _T_23801; // @[LoadQueue.scala 193:43:@8203.6]
  assign _GEN_349 = 3'h7 == _T_23801; // @[LoadQueue.scala 193:43:@8203.6]
  assign _GEN_351 = 3'h1 == _T_23801 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8204.6]
  assign _GEN_352 = 3'h2 == _T_23801 ? shiftedStoreDataKnownPReg_2 : _GEN_351; // @[LoadQueue.scala 194:31:@8204.6]
  assign _GEN_353 = 3'h3 == _T_23801 ? shiftedStoreDataKnownPReg_3 : _GEN_352; // @[LoadQueue.scala 194:31:@8204.6]
  assign _GEN_354 = 3'h4 == _T_23801 ? shiftedStoreDataKnownPReg_4 : _GEN_353; // @[LoadQueue.scala 194:31:@8204.6]
  assign _GEN_355 = 3'h5 == _T_23801 ? shiftedStoreDataKnownPReg_5 : _GEN_354; // @[LoadQueue.scala 194:31:@8204.6]
  assign _GEN_356 = 3'h6 == _T_23801 ? shiftedStoreDataKnownPReg_6 : _GEN_355; // @[LoadQueue.scala 194:31:@8204.6]
  assign _GEN_357 = 3'h7 == _T_23801 ? shiftedStoreDataKnownPReg_7 : _GEN_356; // @[LoadQueue.scala 194:31:@8204.6]
  assign _GEN_359 = 3'h1 == _T_23801 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8205.6]
  assign _GEN_360 = 3'h2 == _T_23801 ? shiftedStoreDataQPreg_2 : _GEN_359; // @[LoadQueue.scala 195:31:@8205.6]
  assign _GEN_361 = 3'h3 == _T_23801 ? shiftedStoreDataQPreg_3 : _GEN_360; // @[LoadQueue.scala 195:31:@8205.6]
  assign _GEN_362 = 3'h4 == _T_23801 ? shiftedStoreDataQPreg_4 : _GEN_361; // @[LoadQueue.scala 195:31:@8205.6]
  assign _GEN_363 = 3'h5 == _T_23801 ? shiftedStoreDataQPreg_5 : _GEN_362; // @[LoadQueue.scala 195:31:@8205.6]
  assign _GEN_364 = 3'h6 == _T_23801 ? shiftedStoreDataQPreg_6 : _GEN_363; // @[LoadQueue.scala 195:31:@8205.6]
  assign _GEN_365 = 3'h7 == _T_23801 ? shiftedStoreDataQPreg_7 : _GEN_364; // @[LoadQueue.scala 195:31:@8205.6]
  assign lastConflict_3_0 = _T_23810 ? _GEN_342 : 1'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign lastConflict_3_1 = _T_23810 ? _GEN_343 : 1'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign lastConflict_3_2 = _T_23810 ? _GEN_344 : 1'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign lastConflict_3_3 = _T_23810 ? _GEN_345 : 1'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign lastConflict_3_4 = _T_23810 ? _GEN_346 : 1'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign lastConflict_3_5 = _T_23810 ? _GEN_347 : 1'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign lastConflict_3_6 = _T_23810 ? _GEN_348 : 1'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign lastConflict_3_7 = _T_23810 ? _GEN_349 : 1'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign canBypass_3 = _T_23810 ? _GEN_357 : 1'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign bypassVal_3 = _T_23810 ? _GEN_365 : 32'h0; // @[LoadQueue.scala 192:53:@8202.4]
  assign _T_23876 = conflictPReg_4_2 ? 2'h2 : {{1'd0}, conflictPReg_4_1}; // @[LoadQueue.scala 191:60:@8235.4]
  assign _T_23877 = conflictPReg_4_3 ? 2'h3 : _T_23876; // @[LoadQueue.scala 191:60:@8236.4]
  assign _T_23878 = conflictPReg_4_4 ? 3'h4 : {{1'd0}, _T_23877}; // @[LoadQueue.scala 191:60:@8237.4]
  assign _T_23879 = conflictPReg_4_5 ? 3'h5 : _T_23878; // @[LoadQueue.scala 191:60:@8238.4]
  assign _T_23880 = conflictPReg_4_6 ? 3'h6 : _T_23879; // @[LoadQueue.scala 191:60:@8239.4]
  assign _T_23881 = conflictPReg_4_7 ? 3'h7 : _T_23880; // @[LoadQueue.scala 191:60:@8240.4]
  assign _T_23884 = conflictPReg_4_0 | conflictPReg_4_1; // @[LoadQueue.scala 192:43:@8242.4]
  assign _T_23885 = _T_23884 | conflictPReg_4_2; // @[LoadQueue.scala 192:43:@8243.4]
  assign _T_23886 = _T_23885 | conflictPReg_4_3; // @[LoadQueue.scala 192:43:@8244.4]
  assign _T_23887 = _T_23886 | conflictPReg_4_4; // @[LoadQueue.scala 192:43:@8245.4]
  assign _T_23888 = _T_23887 | conflictPReg_4_5; // @[LoadQueue.scala 192:43:@8246.4]
  assign _T_23889 = _T_23888 | conflictPReg_4_6; // @[LoadQueue.scala 192:43:@8247.4]
  assign _T_23890 = _T_23889 | conflictPReg_4_7; // @[LoadQueue.scala 192:43:@8248.4]
  assign _GEN_376 = 3'h0 == _T_23881; // @[LoadQueue.scala 193:43:@8250.6]
  assign _GEN_377 = 3'h1 == _T_23881; // @[LoadQueue.scala 193:43:@8250.6]
  assign _GEN_378 = 3'h2 == _T_23881; // @[LoadQueue.scala 193:43:@8250.6]
  assign _GEN_379 = 3'h3 == _T_23881; // @[LoadQueue.scala 193:43:@8250.6]
  assign _GEN_380 = 3'h4 == _T_23881; // @[LoadQueue.scala 193:43:@8250.6]
  assign _GEN_381 = 3'h5 == _T_23881; // @[LoadQueue.scala 193:43:@8250.6]
  assign _GEN_382 = 3'h6 == _T_23881; // @[LoadQueue.scala 193:43:@8250.6]
  assign _GEN_383 = 3'h7 == _T_23881; // @[LoadQueue.scala 193:43:@8250.6]
  assign _GEN_385 = 3'h1 == _T_23881 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8251.6]
  assign _GEN_386 = 3'h2 == _T_23881 ? shiftedStoreDataKnownPReg_2 : _GEN_385; // @[LoadQueue.scala 194:31:@8251.6]
  assign _GEN_387 = 3'h3 == _T_23881 ? shiftedStoreDataKnownPReg_3 : _GEN_386; // @[LoadQueue.scala 194:31:@8251.6]
  assign _GEN_388 = 3'h4 == _T_23881 ? shiftedStoreDataKnownPReg_4 : _GEN_387; // @[LoadQueue.scala 194:31:@8251.6]
  assign _GEN_389 = 3'h5 == _T_23881 ? shiftedStoreDataKnownPReg_5 : _GEN_388; // @[LoadQueue.scala 194:31:@8251.6]
  assign _GEN_390 = 3'h6 == _T_23881 ? shiftedStoreDataKnownPReg_6 : _GEN_389; // @[LoadQueue.scala 194:31:@8251.6]
  assign _GEN_391 = 3'h7 == _T_23881 ? shiftedStoreDataKnownPReg_7 : _GEN_390; // @[LoadQueue.scala 194:31:@8251.6]
  assign _GEN_393 = 3'h1 == _T_23881 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8252.6]
  assign _GEN_394 = 3'h2 == _T_23881 ? shiftedStoreDataQPreg_2 : _GEN_393; // @[LoadQueue.scala 195:31:@8252.6]
  assign _GEN_395 = 3'h3 == _T_23881 ? shiftedStoreDataQPreg_3 : _GEN_394; // @[LoadQueue.scala 195:31:@8252.6]
  assign _GEN_396 = 3'h4 == _T_23881 ? shiftedStoreDataQPreg_4 : _GEN_395; // @[LoadQueue.scala 195:31:@8252.6]
  assign _GEN_397 = 3'h5 == _T_23881 ? shiftedStoreDataQPreg_5 : _GEN_396; // @[LoadQueue.scala 195:31:@8252.6]
  assign _GEN_398 = 3'h6 == _T_23881 ? shiftedStoreDataQPreg_6 : _GEN_397; // @[LoadQueue.scala 195:31:@8252.6]
  assign _GEN_399 = 3'h7 == _T_23881 ? shiftedStoreDataQPreg_7 : _GEN_398; // @[LoadQueue.scala 195:31:@8252.6]
  assign lastConflict_4_0 = _T_23890 ? _GEN_376 : 1'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign lastConflict_4_1 = _T_23890 ? _GEN_377 : 1'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign lastConflict_4_2 = _T_23890 ? _GEN_378 : 1'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign lastConflict_4_3 = _T_23890 ? _GEN_379 : 1'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign lastConflict_4_4 = _T_23890 ? _GEN_380 : 1'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign lastConflict_4_5 = _T_23890 ? _GEN_381 : 1'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign lastConflict_4_6 = _T_23890 ? _GEN_382 : 1'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign lastConflict_4_7 = _T_23890 ? _GEN_383 : 1'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign canBypass_4 = _T_23890 ? _GEN_391 : 1'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign bypassVal_4 = _T_23890 ? _GEN_399 : 32'h0; // @[LoadQueue.scala 192:53:@8249.4]
  assign _T_23956 = conflictPReg_5_2 ? 2'h2 : {{1'd0}, conflictPReg_5_1}; // @[LoadQueue.scala 191:60:@8282.4]
  assign _T_23957 = conflictPReg_5_3 ? 2'h3 : _T_23956; // @[LoadQueue.scala 191:60:@8283.4]
  assign _T_23958 = conflictPReg_5_4 ? 3'h4 : {{1'd0}, _T_23957}; // @[LoadQueue.scala 191:60:@8284.4]
  assign _T_23959 = conflictPReg_5_5 ? 3'h5 : _T_23958; // @[LoadQueue.scala 191:60:@8285.4]
  assign _T_23960 = conflictPReg_5_6 ? 3'h6 : _T_23959; // @[LoadQueue.scala 191:60:@8286.4]
  assign _T_23961 = conflictPReg_5_7 ? 3'h7 : _T_23960; // @[LoadQueue.scala 191:60:@8287.4]
  assign _T_23964 = conflictPReg_5_0 | conflictPReg_5_1; // @[LoadQueue.scala 192:43:@8289.4]
  assign _T_23965 = _T_23964 | conflictPReg_5_2; // @[LoadQueue.scala 192:43:@8290.4]
  assign _T_23966 = _T_23965 | conflictPReg_5_3; // @[LoadQueue.scala 192:43:@8291.4]
  assign _T_23967 = _T_23966 | conflictPReg_5_4; // @[LoadQueue.scala 192:43:@8292.4]
  assign _T_23968 = _T_23967 | conflictPReg_5_5; // @[LoadQueue.scala 192:43:@8293.4]
  assign _T_23969 = _T_23968 | conflictPReg_5_6; // @[LoadQueue.scala 192:43:@8294.4]
  assign _T_23970 = _T_23969 | conflictPReg_5_7; // @[LoadQueue.scala 192:43:@8295.4]
  assign _GEN_410 = 3'h0 == _T_23961; // @[LoadQueue.scala 193:43:@8297.6]
  assign _GEN_411 = 3'h1 == _T_23961; // @[LoadQueue.scala 193:43:@8297.6]
  assign _GEN_412 = 3'h2 == _T_23961; // @[LoadQueue.scala 193:43:@8297.6]
  assign _GEN_413 = 3'h3 == _T_23961; // @[LoadQueue.scala 193:43:@8297.6]
  assign _GEN_414 = 3'h4 == _T_23961; // @[LoadQueue.scala 193:43:@8297.6]
  assign _GEN_415 = 3'h5 == _T_23961; // @[LoadQueue.scala 193:43:@8297.6]
  assign _GEN_416 = 3'h6 == _T_23961; // @[LoadQueue.scala 193:43:@8297.6]
  assign _GEN_417 = 3'h7 == _T_23961; // @[LoadQueue.scala 193:43:@8297.6]
  assign _GEN_419 = 3'h1 == _T_23961 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8298.6]
  assign _GEN_420 = 3'h2 == _T_23961 ? shiftedStoreDataKnownPReg_2 : _GEN_419; // @[LoadQueue.scala 194:31:@8298.6]
  assign _GEN_421 = 3'h3 == _T_23961 ? shiftedStoreDataKnownPReg_3 : _GEN_420; // @[LoadQueue.scala 194:31:@8298.6]
  assign _GEN_422 = 3'h4 == _T_23961 ? shiftedStoreDataKnownPReg_4 : _GEN_421; // @[LoadQueue.scala 194:31:@8298.6]
  assign _GEN_423 = 3'h5 == _T_23961 ? shiftedStoreDataKnownPReg_5 : _GEN_422; // @[LoadQueue.scala 194:31:@8298.6]
  assign _GEN_424 = 3'h6 == _T_23961 ? shiftedStoreDataKnownPReg_6 : _GEN_423; // @[LoadQueue.scala 194:31:@8298.6]
  assign _GEN_425 = 3'h7 == _T_23961 ? shiftedStoreDataKnownPReg_7 : _GEN_424; // @[LoadQueue.scala 194:31:@8298.6]
  assign _GEN_427 = 3'h1 == _T_23961 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8299.6]
  assign _GEN_428 = 3'h2 == _T_23961 ? shiftedStoreDataQPreg_2 : _GEN_427; // @[LoadQueue.scala 195:31:@8299.6]
  assign _GEN_429 = 3'h3 == _T_23961 ? shiftedStoreDataQPreg_3 : _GEN_428; // @[LoadQueue.scala 195:31:@8299.6]
  assign _GEN_430 = 3'h4 == _T_23961 ? shiftedStoreDataQPreg_4 : _GEN_429; // @[LoadQueue.scala 195:31:@8299.6]
  assign _GEN_431 = 3'h5 == _T_23961 ? shiftedStoreDataQPreg_5 : _GEN_430; // @[LoadQueue.scala 195:31:@8299.6]
  assign _GEN_432 = 3'h6 == _T_23961 ? shiftedStoreDataQPreg_6 : _GEN_431; // @[LoadQueue.scala 195:31:@8299.6]
  assign _GEN_433 = 3'h7 == _T_23961 ? shiftedStoreDataQPreg_7 : _GEN_432; // @[LoadQueue.scala 195:31:@8299.6]
  assign lastConflict_5_0 = _T_23970 ? _GEN_410 : 1'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign lastConflict_5_1 = _T_23970 ? _GEN_411 : 1'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign lastConflict_5_2 = _T_23970 ? _GEN_412 : 1'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign lastConflict_5_3 = _T_23970 ? _GEN_413 : 1'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign lastConflict_5_4 = _T_23970 ? _GEN_414 : 1'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign lastConflict_5_5 = _T_23970 ? _GEN_415 : 1'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign lastConflict_5_6 = _T_23970 ? _GEN_416 : 1'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign lastConflict_5_7 = _T_23970 ? _GEN_417 : 1'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign canBypass_5 = _T_23970 ? _GEN_425 : 1'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign bypassVal_5 = _T_23970 ? _GEN_433 : 32'h0; // @[LoadQueue.scala 192:53:@8296.4]
  assign _T_24036 = conflictPReg_6_2 ? 2'h2 : {{1'd0}, conflictPReg_6_1}; // @[LoadQueue.scala 191:60:@8329.4]
  assign _T_24037 = conflictPReg_6_3 ? 2'h3 : _T_24036; // @[LoadQueue.scala 191:60:@8330.4]
  assign _T_24038 = conflictPReg_6_4 ? 3'h4 : {{1'd0}, _T_24037}; // @[LoadQueue.scala 191:60:@8331.4]
  assign _T_24039 = conflictPReg_6_5 ? 3'h5 : _T_24038; // @[LoadQueue.scala 191:60:@8332.4]
  assign _T_24040 = conflictPReg_6_6 ? 3'h6 : _T_24039; // @[LoadQueue.scala 191:60:@8333.4]
  assign _T_24041 = conflictPReg_6_7 ? 3'h7 : _T_24040; // @[LoadQueue.scala 191:60:@8334.4]
  assign _T_24044 = conflictPReg_6_0 | conflictPReg_6_1; // @[LoadQueue.scala 192:43:@8336.4]
  assign _T_24045 = _T_24044 | conflictPReg_6_2; // @[LoadQueue.scala 192:43:@8337.4]
  assign _T_24046 = _T_24045 | conflictPReg_6_3; // @[LoadQueue.scala 192:43:@8338.4]
  assign _T_24047 = _T_24046 | conflictPReg_6_4; // @[LoadQueue.scala 192:43:@8339.4]
  assign _T_24048 = _T_24047 | conflictPReg_6_5; // @[LoadQueue.scala 192:43:@8340.4]
  assign _T_24049 = _T_24048 | conflictPReg_6_6; // @[LoadQueue.scala 192:43:@8341.4]
  assign _T_24050 = _T_24049 | conflictPReg_6_7; // @[LoadQueue.scala 192:43:@8342.4]
  assign _GEN_444 = 3'h0 == _T_24041; // @[LoadQueue.scala 193:43:@8344.6]
  assign _GEN_445 = 3'h1 == _T_24041; // @[LoadQueue.scala 193:43:@8344.6]
  assign _GEN_446 = 3'h2 == _T_24041; // @[LoadQueue.scala 193:43:@8344.6]
  assign _GEN_447 = 3'h3 == _T_24041; // @[LoadQueue.scala 193:43:@8344.6]
  assign _GEN_448 = 3'h4 == _T_24041; // @[LoadQueue.scala 193:43:@8344.6]
  assign _GEN_449 = 3'h5 == _T_24041; // @[LoadQueue.scala 193:43:@8344.6]
  assign _GEN_450 = 3'h6 == _T_24041; // @[LoadQueue.scala 193:43:@8344.6]
  assign _GEN_451 = 3'h7 == _T_24041; // @[LoadQueue.scala 193:43:@8344.6]
  assign _GEN_453 = 3'h1 == _T_24041 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8345.6]
  assign _GEN_454 = 3'h2 == _T_24041 ? shiftedStoreDataKnownPReg_2 : _GEN_453; // @[LoadQueue.scala 194:31:@8345.6]
  assign _GEN_455 = 3'h3 == _T_24041 ? shiftedStoreDataKnownPReg_3 : _GEN_454; // @[LoadQueue.scala 194:31:@8345.6]
  assign _GEN_456 = 3'h4 == _T_24041 ? shiftedStoreDataKnownPReg_4 : _GEN_455; // @[LoadQueue.scala 194:31:@8345.6]
  assign _GEN_457 = 3'h5 == _T_24041 ? shiftedStoreDataKnownPReg_5 : _GEN_456; // @[LoadQueue.scala 194:31:@8345.6]
  assign _GEN_458 = 3'h6 == _T_24041 ? shiftedStoreDataKnownPReg_6 : _GEN_457; // @[LoadQueue.scala 194:31:@8345.6]
  assign _GEN_459 = 3'h7 == _T_24041 ? shiftedStoreDataKnownPReg_7 : _GEN_458; // @[LoadQueue.scala 194:31:@8345.6]
  assign _GEN_461 = 3'h1 == _T_24041 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8346.6]
  assign _GEN_462 = 3'h2 == _T_24041 ? shiftedStoreDataQPreg_2 : _GEN_461; // @[LoadQueue.scala 195:31:@8346.6]
  assign _GEN_463 = 3'h3 == _T_24041 ? shiftedStoreDataQPreg_3 : _GEN_462; // @[LoadQueue.scala 195:31:@8346.6]
  assign _GEN_464 = 3'h4 == _T_24041 ? shiftedStoreDataQPreg_4 : _GEN_463; // @[LoadQueue.scala 195:31:@8346.6]
  assign _GEN_465 = 3'h5 == _T_24041 ? shiftedStoreDataQPreg_5 : _GEN_464; // @[LoadQueue.scala 195:31:@8346.6]
  assign _GEN_466 = 3'h6 == _T_24041 ? shiftedStoreDataQPreg_6 : _GEN_465; // @[LoadQueue.scala 195:31:@8346.6]
  assign _GEN_467 = 3'h7 == _T_24041 ? shiftedStoreDataQPreg_7 : _GEN_466; // @[LoadQueue.scala 195:31:@8346.6]
  assign lastConflict_6_0 = _T_24050 ? _GEN_444 : 1'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign lastConflict_6_1 = _T_24050 ? _GEN_445 : 1'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign lastConflict_6_2 = _T_24050 ? _GEN_446 : 1'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign lastConflict_6_3 = _T_24050 ? _GEN_447 : 1'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign lastConflict_6_4 = _T_24050 ? _GEN_448 : 1'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign lastConflict_6_5 = _T_24050 ? _GEN_449 : 1'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign lastConflict_6_6 = _T_24050 ? _GEN_450 : 1'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign lastConflict_6_7 = _T_24050 ? _GEN_451 : 1'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign canBypass_6 = _T_24050 ? _GEN_459 : 1'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign bypassVal_6 = _T_24050 ? _GEN_467 : 32'h0; // @[LoadQueue.scala 192:53:@8343.4]
  assign _T_24116 = conflictPReg_7_2 ? 2'h2 : {{1'd0}, conflictPReg_7_1}; // @[LoadQueue.scala 191:60:@8376.4]
  assign _T_24117 = conflictPReg_7_3 ? 2'h3 : _T_24116; // @[LoadQueue.scala 191:60:@8377.4]
  assign _T_24118 = conflictPReg_7_4 ? 3'h4 : {{1'd0}, _T_24117}; // @[LoadQueue.scala 191:60:@8378.4]
  assign _T_24119 = conflictPReg_7_5 ? 3'h5 : _T_24118; // @[LoadQueue.scala 191:60:@8379.4]
  assign _T_24120 = conflictPReg_7_6 ? 3'h6 : _T_24119; // @[LoadQueue.scala 191:60:@8380.4]
  assign _T_24121 = conflictPReg_7_7 ? 3'h7 : _T_24120; // @[LoadQueue.scala 191:60:@8381.4]
  assign _T_24124 = conflictPReg_7_0 | conflictPReg_7_1; // @[LoadQueue.scala 192:43:@8383.4]
  assign _T_24125 = _T_24124 | conflictPReg_7_2; // @[LoadQueue.scala 192:43:@8384.4]
  assign _T_24126 = _T_24125 | conflictPReg_7_3; // @[LoadQueue.scala 192:43:@8385.4]
  assign _T_24127 = _T_24126 | conflictPReg_7_4; // @[LoadQueue.scala 192:43:@8386.4]
  assign _T_24128 = _T_24127 | conflictPReg_7_5; // @[LoadQueue.scala 192:43:@8387.4]
  assign _T_24129 = _T_24128 | conflictPReg_7_6; // @[LoadQueue.scala 192:43:@8388.4]
  assign _T_24130 = _T_24129 | conflictPReg_7_7; // @[LoadQueue.scala 192:43:@8389.4]
  assign _GEN_478 = 3'h0 == _T_24121; // @[LoadQueue.scala 193:43:@8391.6]
  assign _GEN_479 = 3'h1 == _T_24121; // @[LoadQueue.scala 193:43:@8391.6]
  assign _GEN_480 = 3'h2 == _T_24121; // @[LoadQueue.scala 193:43:@8391.6]
  assign _GEN_481 = 3'h3 == _T_24121; // @[LoadQueue.scala 193:43:@8391.6]
  assign _GEN_482 = 3'h4 == _T_24121; // @[LoadQueue.scala 193:43:@8391.6]
  assign _GEN_483 = 3'h5 == _T_24121; // @[LoadQueue.scala 193:43:@8391.6]
  assign _GEN_484 = 3'h6 == _T_24121; // @[LoadQueue.scala 193:43:@8391.6]
  assign _GEN_485 = 3'h7 == _T_24121; // @[LoadQueue.scala 193:43:@8391.6]
  assign _GEN_487 = 3'h1 == _T_24121 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8392.6]
  assign _GEN_488 = 3'h2 == _T_24121 ? shiftedStoreDataKnownPReg_2 : _GEN_487; // @[LoadQueue.scala 194:31:@8392.6]
  assign _GEN_489 = 3'h3 == _T_24121 ? shiftedStoreDataKnownPReg_3 : _GEN_488; // @[LoadQueue.scala 194:31:@8392.6]
  assign _GEN_490 = 3'h4 == _T_24121 ? shiftedStoreDataKnownPReg_4 : _GEN_489; // @[LoadQueue.scala 194:31:@8392.6]
  assign _GEN_491 = 3'h5 == _T_24121 ? shiftedStoreDataKnownPReg_5 : _GEN_490; // @[LoadQueue.scala 194:31:@8392.6]
  assign _GEN_492 = 3'h6 == _T_24121 ? shiftedStoreDataKnownPReg_6 : _GEN_491; // @[LoadQueue.scala 194:31:@8392.6]
  assign _GEN_493 = 3'h7 == _T_24121 ? shiftedStoreDataKnownPReg_7 : _GEN_492; // @[LoadQueue.scala 194:31:@8392.6]
  assign _GEN_495 = 3'h1 == _T_24121 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8393.6]
  assign _GEN_496 = 3'h2 == _T_24121 ? shiftedStoreDataQPreg_2 : _GEN_495; // @[LoadQueue.scala 195:31:@8393.6]
  assign _GEN_497 = 3'h3 == _T_24121 ? shiftedStoreDataQPreg_3 : _GEN_496; // @[LoadQueue.scala 195:31:@8393.6]
  assign _GEN_498 = 3'h4 == _T_24121 ? shiftedStoreDataQPreg_4 : _GEN_497; // @[LoadQueue.scala 195:31:@8393.6]
  assign _GEN_499 = 3'h5 == _T_24121 ? shiftedStoreDataQPreg_5 : _GEN_498; // @[LoadQueue.scala 195:31:@8393.6]
  assign _GEN_500 = 3'h6 == _T_24121 ? shiftedStoreDataQPreg_6 : _GEN_499; // @[LoadQueue.scala 195:31:@8393.6]
  assign _GEN_501 = 3'h7 == _T_24121 ? shiftedStoreDataQPreg_7 : _GEN_500; // @[LoadQueue.scala 195:31:@8393.6]
  assign lastConflict_7_0 = _T_24130 ? _GEN_478 : 1'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign lastConflict_7_1 = _T_24130 ? _GEN_479 : 1'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign lastConflict_7_2 = _T_24130 ? _GEN_480 : 1'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign lastConflict_7_3 = _T_24130 ? _GEN_481 : 1'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign lastConflict_7_4 = _T_24130 ? _GEN_482 : 1'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign lastConflict_7_5 = _T_24130 ? _GEN_483 : 1'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign lastConflict_7_6 = _T_24130 ? _GEN_484 : 1'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign lastConflict_7_7 = _T_24130 ? _GEN_485 : 1'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign canBypass_7 = _T_24130 ? _GEN_493 : 1'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign bypassVal_7 = _T_24130 ? _GEN_501 : 32'h0; // @[LoadQueue.scala 192:53:@8390.4]
  assign _T_24174 = 8'h1 << head; // @[OneHot.scala 52:12:@8398.4]
  assign _T_24176 = _T_24174[0]; // @[util.scala 33:60:@8400.4]
  assign _T_24177 = _T_24174[1]; // @[util.scala 33:60:@8401.4]
  assign _T_24178 = _T_24174[2]; // @[util.scala 33:60:@8402.4]
  assign _T_24179 = _T_24174[3]; // @[util.scala 33:60:@8403.4]
  assign _T_24180 = _T_24174[4]; // @[util.scala 33:60:@8404.4]
  assign _T_24181 = _T_24174[5]; // @[util.scala 33:60:@8405.4]
  assign _T_24182 = _T_24174[6]; // @[util.scala 33:60:@8406.4]
  assign _T_24183 = _T_24174[7]; // @[util.scala 33:60:@8407.4]
  assign _T_25168 = dataKnownPReg_7 == 1'h0; // @[LoadQueue.scala 229:41:@9154.4]
  assign _T_25169 = addrKnownPReg_7 & _T_25168; // @[LoadQueue.scala 229:38:@9155.4]
  assign _T_25171 = bypassInitiated_7 == 1'h0; // @[LoadQueue.scala 230:12:@9157.6]
  assign _T_25173 = prevPriorityRequest_7 == 1'h0; // @[LoadQueue.scala 230:46:@9158.6]
  assign _T_25174 = _T_25171 & _T_25173; // @[LoadQueue.scala 230:43:@9159.6]
  assign _T_25176 = dataKnown_7 == 1'h0; // @[LoadQueue.scala 230:84:@9160.6]
  assign _T_25177 = _T_25174 & _T_25176; // @[LoadQueue.scala 230:81:@9161.6]
  assign _T_25180 = storeAddrNotKnownFlagsPReg_7_0 | storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 233:86:@9164.8]
  assign _T_25181 = _T_25180 | storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 233:86:@9165.8]
  assign _T_25182 = _T_25181 | storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 233:86:@9166.8]
  assign _T_25183 = _T_25182 | storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 233:86:@9167.8]
  assign _T_25184 = _T_25183 | storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 233:86:@9168.8]
  assign _T_25185 = _T_25184 | storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 233:86:@9169.8]
  assign _T_25186 = _T_25185 | storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 233:86:@9170.8]
  assign _T_25188 = _T_25186 == 1'h0; // @[LoadQueue.scala 233:38:@9171.8]
  assign _T_25199 = _T_24130 == 1'h0; // @[LoadQueue.scala 234:11:@9180.8]
  assign _T_25200 = _T_25188 & _T_25199; // @[LoadQueue.scala 233:103:@9181.8]
  assign _GEN_564 = _T_25177 ? _T_25200 : 1'h0; // @[LoadQueue.scala 230:110:@9162.6]
  assign loadRequest_7 = _T_25169 ? _GEN_564 : 1'h0; // @[LoadQueue.scala 229:71:@9156.4]
  assign _T_24208 = loadRequest_7 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@8417.4]
  assign _T_25116 = dataKnownPReg_6 == 1'h0; // @[LoadQueue.scala 229:41:@9104.4]
  assign _T_25117 = addrKnownPReg_6 & _T_25116; // @[LoadQueue.scala 229:38:@9105.4]
  assign _T_25119 = bypassInitiated_6 == 1'h0; // @[LoadQueue.scala 230:12:@9107.6]
  assign _T_25121 = prevPriorityRequest_6 == 1'h0; // @[LoadQueue.scala 230:46:@9108.6]
  assign _T_25122 = _T_25119 & _T_25121; // @[LoadQueue.scala 230:43:@9109.6]
  assign _T_25124 = dataKnown_6 == 1'h0; // @[LoadQueue.scala 230:84:@9110.6]
  assign _T_25125 = _T_25122 & _T_25124; // @[LoadQueue.scala 230:81:@9111.6]
  assign _T_25128 = storeAddrNotKnownFlagsPReg_6_0 | storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 233:86:@9114.8]
  assign _T_25129 = _T_25128 | storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 233:86:@9115.8]
  assign _T_25130 = _T_25129 | storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 233:86:@9116.8]
  assign _T_25131 = _T_25130 | storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 233:86:@9117.8]
  assign _T_25132 = _T_25131 | storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 233:86:@9118.8]
  assign _T_25133 = _T_25132 | storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 233:86:@9119.8]
  assign _T_25134 = _T_25133 | storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 233:86:@9120.8]
  assign _T_25136 = _T_25134 == 1'h0; // @[LoadQueue.scala 233:38:@9121.8]
  assign _T_25147 = _T_24050 == 1'h0; // @[LoadQueue.scala 234:11:@9130.8]
  assign _T_25148 = _T_25136 & _T_25147; // @[LoadQueue.scala 233:103:@9131.8]
  assign _GEN_560 = _T_25125 ? _T_25148 : 1'h0; // @[LoadQueue.scala 230:110:@9112.6]
  assign loadRequest_6 = _T_25117 ? _GEN_560 : 1'h0; // @[LoadQueue.scala 229:71:@9106.4]
  assign _T_24209 = loadRequest_6 ? 8'h40 : _T_24208; // @[Mux.scala 31:69:@8418.4]
  assign _T_25064 = dataKnownPReg_5 == 1'h0; // @[LoadQueue.scala 229:41:@9054.4]
  assign _T_25065 = addrKnownPReg_5 & _T_25064; // @[LoadQueue.scala 229:38:@9055.4]
  assign _T_25067 = bypassInitiated_5 == 1'h0; // @[LoadQueue.scala 230:12:@9057.6]
  assign _T_25069 = prevPriorityRequest_5 == 1'h0; // @[LoadQueue.scala 230:46:@9058.6]
  assign _T_25070 = _T_25067 & _T_25069; // @[LoadQueue.scala 230:43:@9059.6]
  assign _T_25072 = dataKnown_5 == 1'h0; // @[LoadQueue.scala 230:84:@9060.6]
  assign _T_25073 = _T_25070 & _T_25072; // @[LoadQueue.scala 230:81:@9061.6]
  assign _T_25076 = storeAddrNotKnownFlagsPReg_5_0 | storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 233:86:@9064.8]
  assign _T_25077 = _T_25076 | storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 233:86:@9065.8]
  assign _T_25078 = _T_25077 | storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 233:86:@9066.8]
  assign _T_25079 = _T_25078 | storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 233:86:@9067.8]
  assign _T_25080 = _T_25079 | storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 233:86:@9068.8]
  assign _T_25081 = _T_25080 | storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 233:86:@9069.8]
  assign _T_25082 = _T_25081 | storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 233:86:@9070.8]
  assign _T_25084 = _T_25082 == 1'h0; // @[LoadQueue.scala 233:38:@9071.8]
  assign _T_25095 = _T_23970 == 1'h0; // @[LoadQueue.scala 234:11:@9080.8]
  assign _T_25096 = _T_25084 & _T_25095; // @[LoadQueue.scala 233:103:@9081.8]
  assign _GEN_556 = _T_25073 ? _T_25096 : 1'h0; // @[LoadQueue.scala 230:110:@9062.6]
  assign loadRequest_5 = _T_25065 ? _GEN_556 : 1'h0; // @[LoadQueue.scala 229:71:@9056.4]
  assign _T_24210 = loadRequest_5 ? 8'h20 : _T_24209; // @[Mux.scala 31:69:@8419.4]
  assign _T_25012 = dataKnownPReg_4 == 1'h0; // @[LoadQueue.scala 229:41:@9004.4]
  assign _T_25013 = addrKnownPReg_4 & _T_25012; // @[LoadQueue.scala 229:38:@9005.4]
  assign _T_25015 = bypassInitiated_4 == 1'h0; // @[LoadQueue.scala 230:12:@9007.6]
  assign _T_25017 = prevPriorityRequest_4 == 1'h0; // @[LoadQueue.scala 230:46:@9008.6]
  assign _T_25018 = _T_25015 & _T_25017; // @[LoadQueue.scala 230:43:@9009.6]
  assign _T_25020 = dataKnown_4 == 1'h0; // @[LoadQueue.scala 230:84:@9010.6]
  assign _T_25021 = _T_25018 & _T_25020; // @[LoadQueue.scala 230:81:@9011.6]
  assign _T_25024 = storeAddrNotKnownFlagsPReg_4_0 | storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 233:86:@9014.8]
  assign _T_25025 = _T_25024 | storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 233:86:@9015.8]
  assign _T_25026 = _T_25025 | storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 233:86:@9016.8]
  assign _T_25027 = _T_25026 | storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 233:86:@9017.8]
  assign _T_25028 = _T_25027 | storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 233:86:@9018.8]
  assign _T_25029 = _T_25028 | storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 233:86:@9019.8]
  assign _T_25030 = _T_25029 | storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 233:86:@9020.8]
  assign _T_25032 = _T_25030 == 1'h0; // @[LoadQueue.scala 233:38:@9021.8]
  assign _T_25043 = _T_23890 == 1'h0; // @[LoadQueue.scala 234:11:@9030.8]
  assign _T_25044 = _T_25032 & _T_25043; // @[LoadQueue.scala 233:103:@9031.8]
  assign _GEN_552 = _T_25021 ? _T_25044 : 1'h0; // @[LoadQueue.scala 230:110:@9012.6]
  assign loadRequest_4 = _T_25013 ? _GEN_552 : 1'h0; // @[LoadQueue.scala 229:71:@9006.4]
  assign _T_24211 = loadRequest_4 ? 8'h10 : _T_24210; // @[Mux.scala 31:69:@8420.4]
  assign _T_24960 = dataKnownPReg_3 == 1'h0; // @[LoadQueue.scala 229:41:@8954.4]
  assign _T_24961 = addrKnownPReg_3 & _T_24960; // @[LoadQueue.scala 229:38:@8955.4]
  assign _T_24963 = bypassInitiated_3 == 1'h0; // @[LoadQueue.scala 230:12:@8957.6]
  assign _T_24965 = prevPriorityRequest_3 == 1'h0; // @[LoadQueue.scala 230:46:@8958.6]
  assign _T_24966 = _T_24963 & _T_24965; // @[LoadQueue.scala 230:43:@8959.6]
  assign _T_24968 = dataKnown_3 == 1'h0; // @[LoadQueue.scala 230:84:@8960.6]
  assign _T_24969 = _T_24966 & _T_24968; // @[LoadQueue.scala 230:81:@8961.6]
  assign _T_24972 = storeAddrNotKnownFlagsPReg_3_0 | storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 233:86:@8964.8]
  assign _T_24973 = _T_24972 | storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 233:86:@8965.8]
  assign _T_24974 = _T_24973 | storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 233:86:@8966.8]
  assign _T_24975 = _T_24974 | storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 233:86:@8967.8]
  assign _T_24976 = _T_24975 | storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 233:86:@8968.8]
  assign _T_24977 = _T_24976 | storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 233:86:@8969.8]
  assign _T_24978 = _T_24977 | storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 233:86:@8970.8]
  assign _T_24980 = _T_24978 == 1'h0; // @[LoadQueue.scala 233:38:@8971.8]
  assign _T_24991 = _T_23810 == 1'h0; // @[LoadQueue.scala 234:11:@8980.8]
  assign _T_24992 = _T_24980 & _T_24991; // @[LoadQueue.scala 233:103:@8981.8]
  assign _GEN_548 = _T_24969 ? _T_24992 : 1'h0; // @[LoadQueue.scala 230:110:@8962.6]
  assign loadRequest_3 = _T_24961 ? _GEN_548 : 1'h0; // @[LoadQueue.scala 229:71:@8956.4]
  assign _T_24212 = loadRequest_3 ? 8'h8 : _T_24211; // @[Mux.scala 31:69:@8421.4]
  assign _T_24908 = dataKnownPReg_2 == 1'h0; // @[LoadQueue.scala 229:41:@8904.4]
  assign _T_24909 = addrKnownPReg_2 & _T_24908; // @[LoadQueue.scala 229:38:@8905.4]
  assign _T_24911 = bypassInitiated_2 == 1'h0; // @[LoadQueue.scala 230:12:@8907.6]
  assign _T_24913 = prevPriorityRequest_2 == 1'h0; // @[LoadQueue.scala 230:46:@8908.6]
  assign _T_24914 = _T_24911 & _T_24913; // @[LoadQueue.scala 230:43:@8909.6]
  assign _T_24916 = dataKnown_2 == 1'h0; // @[LoadQueue.scala 230:84:@8910.6]
  assign _T_24917 = _T_24914 & _T_24916; // @[LoadQueue.scala 230:81:@8911.6]
  assign _T_24920 = storeAddrNotKnownFlagsPReg_2_0 | storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 233:86:@8914.8]
  assign _T_24921 = _T_24920 | storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 233:86:@8915.8]
  assign _T_24922 = _T_24921 | storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 233:86:@8916.8]
  assign _T_24923 = _T_24922 | storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 233:86:@8917.8]
  assign _T_24924 = _T_24923 | storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 233:86:@8918.8]
  assign _T_24925 = _T_24924 | storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 233:86:@8919.8]
  assign _T_24926 = _T_24925 | storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 233:86:@8920.8]
  assign _T_24928 = _T_24926 == 1'h0; // @[LoadQueue.scala 233:38:@8921.8]
  assign _T_24939 = _T_23730 == 1'h0; // @[LoadQueue.scala 234:11:@8930.8]
  assign _T_24940 = _T_24928 & _T_24939; // @[LoadQueue.scala 233:103:@8931.8]
  assign _GEN_544 = _T_24917 ? _T_24940 : 1'h0; // @[LoadQueue.scala 230:110:@8912.6]
  assign loadRequest_2 = _T_24909 ? _GEN_544 : 1'h0; // @[LoadQueue.scala 229:71:@8906.4]
  assign _T_24213 = loadRequest_2 ? 8'h4 : _T_24212; // @[Mux.scala 31:69:@8422.4]
  assign _T_24856 = dataKnownPReg_1 == 1'h0; // @[LoadQueue.scala 229:41:@8854.4]
  assign _T_24857 = addrKnownPReg_1 & _T_24856; // @[LoadQueue.scala 229:38:@8855.4]
  assign _T_24859 = bypassInitiated_1 == 1'h0; // @[LoadQueue.scala 230:12:@8857.6]
  assign _T_24861 = prevPriorityRequest_1 == 1'h0; // @[LoadQueue.scala 230:46:@8858.6]
  assign _T_24862 = _T_24859 & _T_24861; // @[LoadQueue.scala 230:43:@8859.6]
  assign _T_24864 = dataKnown_1 == 1'h0; // @[LoadQueue.scala 230:84:@8860.6]
  assign _T_24865 = _T_24862 & _T_24864; // @[LoadQueue.scala 230:81:@8861.6]
  assign _T_24868 = storeAddrNotKnownFlagsPReg_1_0 | storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 233:86:@8864.8]
  assign _T_24869 = _T_24868 | storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 233:86:@8865.8]
  assign _T_24870 = _T_24869 | storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 233:86:@8866.8]
  assign _T_24871 = _T_24870 | storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 233:86:@8867.8]
  assign _T_24872 = _T_24871 | storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 233:86:@8868.8]
  assign _T_24873 = _T_24872 | storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 233:86:@8869.8]
  assign _T_24874 = _T_24873 | storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 233:86:@8870.8]
  assign _T_24876 = _T_24874 == 1'h0; // @[LoadQueue.scala 233:38:@8871.8]
  assign _T_24887 = _T_23650 == 1'h0; // @[LoadQueue.scala 234:11:@8880.8]
  assign _T_24888 = _T_24876 & _T_24887; // @[LoadQueue.scala 233:103:@8881.8]
  assign _GEN_540 = _T_24865 ? _T_24888 : 1'h0; // @[LoadQueue.scala 230:110:@8862.6]
  assign loadRequest_1 = _T_24857 ? _GEN_540 : 1'h0; // @[LoadQueue.scala 229:71:@8856.4]
  assign _T_24214 = loadRequest_1 ? 8'h2 : _T_24213; // @[Mux.scala 31:69:@8423.4]
  assign _T_24804 = dataKnownPReg_0 == 1'h0; // @[LoadQueue.scala 229:41:@8804.4]
  assign _T_24805 = addrKnownPReg_0 & _T_24804; // @[LoadQueue.scala 229:38:@8805.4]
  assign _T_24807 = bypassInitiated_0 == 1'h0; // @[LoadQueue.scala 230:12:@8807.6]
  assign _T_24809 = prevPriorityRequest_0 == 1'h0; // @[LoadQueue.scala 230:46:@8808.6]
  assign _T_24810 = _T_24807 & _T_24809; // @[LoadQueue.scala 230:43:@8809.6]
  assign _T_24812 = dataKnown_0 == 1'h0; // @[LoadQueue.scala 230:84:@8810.6]
  assign _T_24813 = _T_24810 & _T_24812; // @[LoadQueue.scala 230:81:@8811.6]
  assign _T_24816 = storeAddrNotKnownFlagsPReg_0_0 | storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 233:86:@8814.8]
  assign _T_24817 = _T_24816 | storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 233:86:@8815.8]
  assign _T_24818 = _T_24817 | storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 233:86:@8816.8]
  assign _T_24819 = _T_24818 | storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 233:86:@8817.8]
  assign _T_24820 = _T_24819 | storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 233:86:@8818.8]
  assign _T_24821 = _T_24820 | storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 233:86:@8819.8]
  assign _T_24822 = _T_24821 | storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 233:86:@8820.8]
  assign _T_24824 = _T_24822 == 1'h0; // @[LoadQueue.scala 233:38:@8821.8]
  assign _T_24835 = _T_23570 == 1'h0; // @[LoadQueue.scala 234:11:@8830.8]
  assign _T_24836 = _T_24824 & _T_24835; // @[LoadQueue.scala 233:103:@8831.8]
  assign _GEN_536 = _T_24813 ? _T_24836 : 1'h0; // @[LoadQueue.scala 230:110:@8812.6]
  assign loadRequest_0 = _T_24805 ? _GEN_536 : 1'h0; // @[LoadQueue.scala 229:71:@8806.4]
  assign _T_24215 = loadRequest_0 ? 8'h1 : _T_24214; // @[Mux.scala 31:69:@8424.4]
  assign _T_24216 = _T_24215[0]; // @[OneHot.scala 66:30:@8425.4]
  assign _T_24217 = _T_24215[1]; // @[OneHot.scala 66:30:@8426.4]
  assign _T_24218 = _T_24215[2]; // @[OneHot.scala 66:30:@8427.4]
  assign _T_24219 = _T_24215[3]; // @[OneHot.scala 66:30:@8428.4]
  assign _T_24220 = _T_24215[4]; // @[OneHot.scala 66:30:@8429.4]
  assign _T_24221 = _T_24215[5]; // @[OneHot.scala 66:30:@8430.4]
  assign _T_24222 = _T_24215[6]; // @[OneHot.scala 66:30:@8431.4]
  assign _T_24223 = _T_24215[7]; // @[OneHot.scala 66:30:@8432.4]
  assign _T_24248 = loadRequest_0 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@8442.4]
  assign _T_24249 = loadRequest_7 ? 8'h40 : _T_24248; // @[Mux.scala 31:69:@8443.4]
  assign _T_24250 = loadRequest_6 ? 8'h20 : _T_24249; // @[Mux.scala 31:69:@8444.4]
  assign _T_24251 = loadRequest_5 ? 8'h10 : _T_24250; // @[Mux.scala 31:69:@8445.4]
  assign _T_24252 = loadRequest_4 ? 8'h8 : _T_24251; // @[Mux.scala 31:69:@8446.4]
  assign _T_24253 = loadRequest_3 ? 8'h4 : _T_24252; // @[Mux.scala 31:69:@8447.4]
  assign _T_24254 = loadRequest_2 ? 8'h2 : _T_24253; // @[Mux.scala 31:69:@8448.4]
  assign _T_24255 = loadRequest_1 ? 8'h1 : _T_24254; // @[Mux.scala 31:69:@8449.4]
  assign _T_24256 = _T_24255[0]; // @[OneHot.scala 66:30:@8450.4]
  assign _T_24257 = _T_24255[1]; // @[OneHot.scala 66:30:@8451.4]
  assign _T_24258 = _T_24255[2]; // @[OneHot.scala 66:30:@8452.4]
  assign _T_24259 = _T_24255[3]; // @[OneHot.scala 66:30:@8453.4]
  assign _T_24260 = _T_24255[4]; // @[OneHot.scala 66:30:@8454.4]
  assign _T_24261 = _T_24255[5]; // @[OneHot.scala 66:30:@8455.4]
  assign _T_24262 = _T_24255[6]; // @[OneHot.scala 66:30:@8456.4]
  assign _T_24263 = _T_24255[7]; // @[OneHot.scala 66:30:@8457.4]
  assign _T_24288 = loadRequest_1 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@8467.4]
  assign _T_24289 = loadRequest_0 ? 8'h40 : _T_24288; // @[Mux.scala 31:69:@8468.4]
  assign _T_24290 = loadRequest_7 ? 8'h20 : _T_24289; // @[Mux.scala 31:69:@8469.4]
  assign _T_24291 = loadRequest_6 ? 8'h10 : _T_24290; // @[Mux.scala 31:69:@8470.4]
  assign _T_24292 = loadRequest_5 ? 8'h8 : _T_24291; // @[Mux.scala 31:69:@8471.4]
  assign _T_24293 = loadRequest_4 ? 8'h4 : _T_24292; // @[Mux.scala 31:69:@8472.4]
  assign _T_24294 = loadRequest_3 ? 8'h2 : _T_24293; // @[Mux.scala 31:69:@8473.4]
  assign _T_24295 = loadRequest_2 ? 8'h1 : _T_24294; // @[Mux.scala 31:69:@8474.4]
  assign _T_24296 = _T_24295[0]; // @[OneHot.scala 66:30:@8475.4]
  assign _T_24297 = _T_24295[1]; // @[OneHot.scala 66:30:@8476.4]
  assign _T_24298 = _T_24295[2]; // @[OneHot.scala 66:30:@8477.4]
  assign _T_24299 = _T_24295[3]; // @[OneHot.scala 66:30:@8478.4]
  assign _T_24300 = _T_24295[4]; // @[OneHot.scala 66:30:@8479.4]
  assign _T_24301 = _T_24295[5]; // @[OneHot.scala 66:30:@8480.4]
  assign _T_24302 = _T_24295[6]; // @[OneHot.scala 66:30:@8481.4]
  assign _T_24303 = _T_24295[7]; // @[OneHot.scala 66:30:@8482.4]
  assign _T_24328 = loadRequest_2 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@8492.4]
  assign _T_24329 = loadRequest_1 ? 8'h40 : _T_24328; // @[Mux.scala 31:69:@8493.4]
  assign _T_24330 = loadRequest_0 ? 8'h20 : _T_24329; // @[Mux.scala 31:69:@8494.4]
  assign _T_24331 = loadRequest_7 ? 8'h10 : _T_24330; // @[Mux.scala 31:69:@8495.4]
  assign _T_24332 = loadRequest_6 ? 8'h8 : _T_24331; // @[Mux.scala 31:69:@8496.4]
  assign _T_24333 = loadRequest_5 ? 8'h4 : _T_24332; // @[Mux.scala 31:69:@8497.4]
  assign _T_24334 = loadRequest_4 ? 8'h2 : _T_24333; // @[Mux.scala 31:69:@8498.4]
  assign _T_24335 = loadRequest_3 ? 8'h1 : _T_24334; // @[Mux.scala 31:69:@8499.4]
  assign _T_24336 = _T_24335[0]; // @[OneHot.scala 66:30:@8500.4]
  assign _T_24337 = _T_24335[1]; // @[OneHot.scala 66:30:@8501.4]
  assign _T_24338 = _T_24335[2]; // @[OneHot.scala 66:30:@8502.4]
  assign _T_24339 = _T_24335[3]; // @[OneHot.scala 66:30:@8503.4]
  assign _T_24340 = _T_24335[4]; // @[OneHot.scala 66:30:@8504.4]
  assign _T_24341 = _T_24335[5]; // @[OneHot.scala 66:30:@8505.4]
  assign _T_24342 = _T_24335[6]; // @[OneHot.scala 66:30:@8506.4]
  assign _T_24343 = _T_24335[7]; // @[OneHot.scala 66:30:@8507.4]
  assign _T_24368 = loadRequest_3 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@8517.4]
  assign _T_24369 = loadRequest_2 ? 8'h40 : _T_24368; // @[Mux.scala 31:69:@8518.4]
  assign _T_24370 = loadRequest_1 ? 8'h20 : _T_24369; // @[Mux.scala 31:69:@8519.4]
  assign _T_24371 = loadRequest_0 ? 8'h10 : _T_24370; // @[Mux.scala 31:69:@8520.4]
  assign _T_24372 = loadRequest_7 ? 8'h8 : _T_24371; // @[Mux.scala 31:69:@8521.4]
  assign _T_24373 = loadRequest_6 ? 8'h4 : _T_24372; // @[Mux.scala 31:69:@8522.4]
  assign _T_24374 = loadRequest_5 ? 8'h2 : _T_24373; // @[Mux.scala 31:69:@8523.4]
  assign _T_24375 = loadRequest_4 ? 8'h1 : _T_24374; // @[Mux.scala 31:69:@8524.4]
  assign _T_24376 = _T_24375[0]; // @[OneHot.scala 66:30:@8525.4]
  assign _T_24377 = _T_24375[1]; // @[OneHot.scala 66:30:@8526.4]
  assign _T_24378 = _T_24375[2]; // @[OneHot.scala 66:30:@8527.4]
  assign _T_24379 = _T_24375[3]; // @[OneHot.scala 66:30:@8528.4]
  assign _T_24380 = _T_24375[4]; // @[OneHot.scala 66:30:@8529.4]
  assign _T_24381 = _T_24375[5]; // @[OneHot.scala 66:30:@8530.4]
  assign _T_24382 = _T_24375[6]; // @[OneHot.scala 66:30:@8531.4]
  assign _T_24383 = _T_24375[7]; // @[OneHot.scala 66:30:@8532.4]
  assign _T_24408 = loadRequest_4 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@8542.4]
  assign _T_24409 = loadRequest_3 ? 8'h40 : _T_24408; // @[Mux.scala 31:69:@8543.4]
  assign _T_24410 = loadRequest_2 ? 8'h20 : _T_24409; // @[Mux.scala 31:69:@8544.4]
  assign _T_24411 = loadRequest_1 ? 8'h10 : _T_24410; // @[Mux.scala 31:69:@8545.4]
  assign _T_24412 = loadRequest_0 ? 8'h8 : _T_24411; // @[Mux.scala 31:69:@8546.4]
  assign _T_24413 = loadRequest_7 ? 8'h4 : _T_24412; // @[Mux.scala 31:69:@8547.4]
  assign _T_24414 = loadRequest_6 ? 8'h2 : _T_24413; // @[Mux.scala 31:69:@8548.4]
  assign _T_24415 = loadRequest_5 ? 8'h1 : _T_24414; // @[Mux.scala 31:69:@8549.4]
  assign _T_24416 = _T_24415[0]; // @[OneHot.scala 66:30:@8550.4]
  assign _T_24417 = _T_24415[1]; // @[OneHot.scala 66:30:@8551.4]
  assign _T_24418 = _T_24415[2]; // @[OneHot.scala 66:30:@8552.4]
  assign _T_24419 = _T_24415[3]; // @[OneHot.scala 66:30:@8553.4]
  assign _T_24420 = _T_24415[4]; // @[OneHot.scala 66:30:@8554.4]
  assign _T_24421 = _T_24415[5]; // @[OneHot.scala 66:30:@8555.4]
  assign _T_24422 = _T_24415[6]; // @[OneHot.scala 66:30:@8556.4]
  assign _T_24423 = _T_24415[7]; // @[OneHot.scala 66:30:@8557.4]
  assign _T_24448 = loadRequest_5 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@8567.4]
  assign _T_24449 = loadRequest_4 ? 8'h40 : _T_24448; // @[Mux.scala 31:69:@8568.4]
  assign _T_24450 = loadRequest_3 ? 8'h20 : _T_24449; // @[Mux.scala 31:69:@8569.4]
  assign _T_24451 = loadRequest_2 ? 8'h10 : _T_24450; // @[Mux.scala 31:69:@8570.4]
  assign _T_24452 = loadRequest_1 ? 8'h8 : _T_24451; // @[Mux.scala 31:69:@8571.4]
  assign _T_24453 = loadRequest_0 ? 8'h4 : _T_24452; // @[Mux.scala 31:69:@8572.4]
  assign _T_24454 = loadRequest_7 ? 8'h2 : _T_24453; // @[Mux.scala 31:69:@8573.4]
  assign _T_24455 = loadRequest_6 ? 8'h1 : _T_24454; // @[Mux.scala 31:69:@8574.4]
  assign _T_24456 = _T_24455[0]; // @[OneHot.scala 66:30:@8575.4]
  assign _T_24457 = _T_24455[1]; // @[OneHot.scala 66:30:@8576.4]
  assign _T_24458 = _T_24455[2]; // @[OneHot.scala 66:30:@8577.4]
  assign _T_24459 = _T_24455[3]; // @[OneHot.scala 66:30:@8578.4]
  assign _T_24460 = _T_24455[4]; // @[OneHot.scala 66:30:@8579.4]
  assign _T_24461 = _T_24455[5]; // @[OneHot.scala 66:30:@8580.4]
  assign _T_24462 = _T_24455[6]; // @[OneHot.scala 66:30:@8581.4]
  assign _T_24463 = _T_24455[7]; // @[OneHot.scala 66:30:@8582.4]
  assign _T_24488 = loadRequest_6 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@8592.4]
  assign _T_24489 = loadRequest_5 ? 8'h40 : _T_24488; // @[Mux.scala 31:69:@8593.4]
  assign _T_24490 = loadRequest_4 ? 8'h20 : _T_24489; // @[Mux.scala 31:69:@8594.4]
  assign _T_24491 = loadRequest_3 ? 8'h10 : _T_24490; // @[Mux.scala 31:69:@8595.4]
  assign _T_24492 = loadRequest_2 ? 8'h8 : _T_24491; // @[Mux.scala 31:69:@8596.4]
  assign _T_24493 = loadRequest_1 ? 8'h4 : _T_24492; // @[Mux.scala 31:69:@8597.4]
  assign _T_24494 = loadRequest_0 ? 8'h2 : _T_24493; // @[Mux.scala 31:69:@8598.4]
  assign _T_24495 = loadRequest_7 ? 8'h1 : _T_24494; // @[Mux.scala 31:69:@8599.4]
  assign _T_24496 = _T_24495[0]; // @[OneHot.scala 66:30:@8600.4]
  assign _T_24497 = _T_24495[1]; // @[OneHot.scala 66:30:@8601.4]
  assign _T_24498 = _T_24495[2]; // @[OneHot.scala 66:30:@8602.4]
  assign _T_24499 = _T_24495[3]; // @[OneHot.scala 66:30:@8603.4]
  assign _T_24500 = _T_24495[4]; // @[OneHot.scala 66:30:@8604.4]
  assign _T_24501 = _T_24495[5]; // @[OneHot.scala 66:30:@8605.4]
  assign _T_24502 = _T_24495[6]; // @[OneHot.scala 66:30:@8606.4]
  assign _T_24503 = _T_24495[7]; // @[OneHot.scala 66:30:@8607.4]
  assign _T_24544 = {_T_24223,_T_24222,_T_24221,_T_24220,_T_24219,_T_24218,_T_24217,_T_24216}; // @[Mux.scala 19:72:@8623.4]
  assign _T_24546 = _T_24176 ? _T_24544 : 8'h0; // @[Mux.scala 19:72:@8624.4]
  assign _T_24553 = {_T_24262,_T_24261,_T_24260,_T_24259,_T_24258,_T_24257,_T_24256,_T_24263}; // @[Mux.scala 19:72:@8631.4]
  assign _T_24555 = _T_24177 ? _T_24553 : 8'h0; // @[Mux.scala 19:72:@8632.4]
  assign _T_24562 = {_T_24301,_T_24300,_T_24299,_T_24298,_T_24297,_T_24296,_T_24303,_T_24302}; // @[Mux.scala 19:72:@8639.4]
  assign _T_24564 = _T_24178 ? _T_24562 : 8'h0; // @[Mux.scala 19:72:@8640.4]
  assign _T_24571 = {_T_24340,_T_24339,_T_24338,_T_24337,_T_24336,_T_24343,_T_24342,_T_24341}; // @[Mux.scala 19:72:@8647.4]
  assign _T_24573 = _T_24179 ? _T_24571 : 8'h0; // @[Mux.scala 19:72:@8648.4]
  assign _T_24580 = {_T_24379,_T_24378,_T_24377,_T_24376,_T_24383,_T_24382,_T_24381,_T_24380}; // @[Mux.scala 19:72:@8655.4]
  assign _T_24582 = _T_24180 ? _T_24580 : 8'h0; // @[Mux.scala 19:72:@8656.4]
  assign _T_24589 = {_T_24418,_T_24417,_T_24416,_T_24423,_T_24422,_T_24421,_T_24420,_T_24419}; // @[Mux.scala 19:72:@8663.4]
  assign _T_24591 = _T_24181 ? _T_24589 : 8'h0; // @[Mux.scala 19:72:@8664.4]
  assign _T_24598 = {_T_24457,_T_24456,_T_24463,_T_24462,_T_24461,_T_24460,_T_24459,_T_24458}; // @[Mux.scala 19:72:@8671.4]
  assign _T_24600 = _T_24182 ? _T_24598 : 8'h0; // @[Mux.scala 19:72:@8672.4]
  assign _T_24607 = {_T_24496,_T_24503,_T_24502,_T_24501,_T_24500,_T_24499,_T_24498,_T_24497}; // @[Mux.scala 19:72:@8679.4]
  assign _T_24609 = _T_24183 ? _T_24607 : 8'h0; // @[Mux.scala 19:72:@8680.4]
  assign _T_24610 = _T_24546 | _T_24555; // @[Mux.scala 19:72:@8681.4]
  assign _T_24611 = _T_24610 | _T_24564; // @[Mux.scala 19:72:@8682.4]
  assign _T_24612 = _T_24611 | _T_24573; // @[Mux.scala 19:72:@8683.4]
  assign _T_24613 = _T_24612 | _T_24582; // @[Mux.scala 19:72:@8684.4]
  assign _T_24614 = _T_24613 | _T_24591; // @[Mux.scala 19:72:@8685.4]
  assign _T_24615 = _T_24614 | _T_24600; // @[Mux.scala 19:72:@8686.4]
  assign _T_24616 = _T_24615 | _T_24609; // @[Mux.scala 19:72:@8687.4]
  assign priorityLoadRequest_0 = _T_24616[0]; // @[Mux.scala 19:72:@8691.4]
  assign priorityLoadRequest_1 = _T_24616[1]; // @[Mux.scala 19:72:@8693.4]
  assign priorityLoadRequest_2 = _T_24616[2]; // @[Mux.scala 19:72:@8695.4]
  assign priorityLoadRequest_3 = _T_24616[3]; // @[Mux.scala 19:72:@8697.4]
  assign priorityLoadRequest_4 = _T_24616[4]; // @[Mux.scala 19:72:@8699.4]
  assign priorityLoadRequest_5 = _T_24616[5]; // @[Mux.scala 19:72:@8701.4]
  assign priorityLoadRequest_6 = _T_24616[6]; // @[Mux.scala 19:72:@8703.4]
  assign priorityLoadRequest_7 = _T_24616[7]; // @[Mux.scala 19:72:@8705.4]
  assign _GEN_512 = io_memIsReadyForLoads ? priorityLoadRequest_0 : 1'h0; // @[LoadQueue.scala 208:31:@8717.4]
  assign _GEN_513 = io_memIsReadyForLoads ? priorityLoadRequest_1 : 1'h0; // @[LoadQueue.scala 208:31:@8717.4]
  assign _GEN_514 = io_memIsReadyForLoads ? priorityLoadRequest_2 : 1'h0; // @[LoadQueue.scala 208:31:@8717.4]
  assign _GEN_515 = io_memIsReadyForLoads ? priorityLoadRequest_3 : 1'h0; // @[LoadQueue.scala 208:31:@8717.4]
  assign _GEN_516 = io_memIsReadyForLoads ? priorityLoadRequest_4 : 1'h0; // @[LoadQueue.scala 208:31:@8717.4]
  assign _GEN_517 = io_memIsReadyForLoads ? priorityLoadRequest_5 : 1'h0; // @[LoadQueue.scala 208:31:@8717.4]
  assign _GEN_518 = io_memIsReadyForLoads ? priorityLoadRequest_6 : 1'h0; // @[LoadQueue.scala 208:31:@8717.4]
  assign _GEN_519 = io_memIsReadyForLoads ? priorityLoadRequest_7 : 1'h0; // @[LoadQueue.scala 208:31:@8717.4]
  assign _T_24843 = {storeAddrNotKnownFlagsPReg_0_7,storeAddrNotKnownFlagsPReg_0_6,storeAddrNotKnownFlagsPReg_0_5,storeAddrNotKnownFlagsPReg_0_4,storeAddrNotKnownFlagsPReg_0_3,storeAddrNotKnownFlagsPReg_0_2,storeAddrNotKnownFlagsPReg_0_1,storeAddrNotKnownFlagsPReg_0_0}; // @[LoadQueue.scala 238:58:@8839.8]
  assign _T_24850 = {lastConflict_0_7,lastConflict_0_6,lastConflict_0_5,lastConflict_0_4,lastConflict_0_3,lastConflict_0_2,lastConflict_0_1,lastConflict_0_0}; // @[LoadQueue.scala 238:96:@8846.8]
  assign _T_24851 = _T_24843 < _T_24850; // @[LoadQueue.scala 238:61:@8847.8]
  assign _T_24852 = canBypass_0 & _T_24851; // @[LoadQueue.scala 237:64:@8848.8]
  assign _GEN_537 = _T_24813 ? _T_24852 : 1'h0; // @[LoadQueue.scala 230:110:@8812.6]
  assign bypassRequest_0 = _T_24805 ? _GEN_537 : 1'h0; // @[LoadQueue.scala 229:71:@8806.4]
  assign _GEN_520 = bypassRequest_0 ? 1'h1 : bypassInitiated_0; // @[LoadQueue.scala 217:34:@8750.6]
  assign _GEN_521 = initBits_0 ? 1'h0 : _GEN_520; // @[LoadQueue.scala 215:23:@8746.4]
  assign _T_24895 = {storeAddrNotKnownFlagsPReg_1_7,storeAddrNotKnownFlagsPReg_1_6,storeAddrNotKnownFlagsPReg_1_5,storeAddrNotKnownFlagsPReg_1_4,storeAddrNotKnownFlagsPReg_1_3,storeAddrNotKnownFlagsPReg_1_2,storeAddrNotKnownFlagsPReg_1_1,storeAddrNotKnownFlagsPReg_1_0}; // @[LoadQueue.scala 238:58:@8889.8]
  assign _T_24902 = {lastConflict_1_7,lastConflict_1_6,lastConflict_1_5,lastConflict_1_4,lastConflict_1_3,lastConflict_1_2,lastConflict_1_1,lastConflict_1_0}; // @[LoadQueue.scala 238:96:@8896.8]
  assign _T_24903 = _T_24895 < _T_24902; // @[LoadQueue.scala 238:61:@8897.8]
  assign _T_24904 = canBypass_1 & _T_24903; // @[LoadQueue.scala 237:64:@8898.8]
  assign _GEN_541 = _T_24865 ? _T_24904 : 1'h0; // @[LoadQueue.scala 230:110:@8862.6]
  assign bypassRequest_1 = _T_24857 ? _GEN_541 : 1'h0; // @[LoadQueue.scala 229:71:@8856.4]
  assign _GEN_522 = bypassRequest_1 ? 1'h1 : bypassInitiated_1; // @[LoadQueue.scala 217:34:@8757.6]
  assign _GEN_523 = initBits_1 ? 1'h0 : _GEN_522; // @[LoadQueue.scala 215:23:@8753.4]
  assign _T_24947 = {storeAddrNotKnownFlagsPReg_2_7,storeAddrNotKnownFlagsPReg_2_6,storeAddrNotKnownFlagsPReg_2_5,storeAddrNotKnownFlagsPReg_2_4,storeAddrNotKnownFlagsPReg_2_3,storeAddrNotKnownFlagsPReg_2_2,storeAddrNotKnownFlagsPReg_2_1,storeAddrNotKnownFlagsPReg_2_0}; // @[LoadQueue.scala 238:58:@8939.8]
  assign _T_24954 = {lastConflict_2_7,lastConflict_2_6,lastConflict_2_5,lastConflict_2_4,lastConflict_2_3,lastConflict_2_2,lastConflict_2_1,lastConflict_2_0}; // @[LoadQueue.scala 238:96:@8946.8]
  assign _T_24955 = _T_24947 < _T_24954; // @[LoadQueue.scala 238:61:@8947.8]
  assign _T_24956 = canBypass_2 & _T_24955; // @[LoadQueue.scala 237:64:@8948.8]
  assign _GEN_545 = _T_24917 ? _T_24956 : 1'h0; // @[LoadQueue.scala 230:110:@8912.6]
  assign bypassRequest_2 = _T_24909 ? _GEN_545 : 1'h0; // @[LoadQueue.scala 229:71:@8906.4]
  assign _GEN_524 = bypassRequest_2 ? 1'h1 : bypassInitiated_2; // @[LoadQueue.scala 217:34:@8764.6]
  assign _GEN_525 = initBits_2 ? 1'h0 : _GEN_524; // @[LoadQueue.scala 215:23:@8760.4]
  assign _T_24999 = {storeAddrNotKnownFlagsPReg_3_7,storeAddrNotKnownFlagsPReg_3_6,storeAddrNotKnownFlagsPReg_3_5,storeAddrNotKnownFlagsPReg_3_4,storeAddrNotKnownFlagsPReg_3_3,storeAddrNotKnownFlagsPReg_3_2,storeAddrNotKnownFlagsPReg_3_1,storeAddrNotKnownFlagsPReg_3_0}; // @[LoadQueue.scala 238:58:@8989.8]
  assign _T_25006 = {lastConflict_3_7,lastConflict_3_6,lastConflict_3_5,lastConflict_3_4,lastConflict_3_3,lastConflict_3_2,lastConflict_3_1,lastConflict_3_0}; // @[LoadQueue.scala 238:96:@8996.8]
  assign _T_25007 = _T_24999 < _T_25006; // @[LoadQueue.scala 238:61:@8997.8]
  assign _T_25008 = canBypass_3 & _T_25007; // @[LoadQueue.scala 237:64:@8998.8]
  assign _GEN_549 = _T_24969 ? _T_25008 : 1'h0; // @[LoadQueue.scala 230:110:@8962.6]
  assign bypassRequest_3 = _T_24961 ? _GEN_549 : 1'h0; // @[LoadQueue.scala 229:71:@8956.4]
  assign _GEN_526 = bypassRequest_3 ? 1'h1 : bypassInitiated_3; // @[LoadQueue.scala 217:34:@8771.6]
  assign _GEN_527 = initBits_3 ? 1'h0 : _GEN_526; // @[LoadQueue.scala 215:23:@8767.4]
  assign _T_25051 = {storeAddrNotKnownFlagsPReg_4_7,storeAddrNotKnownFlagsPReg_4_6,storeAddrNotKnownFlagsPReg_4_5,storeAddrNotKnownFlagsPReg_4_4,storeAddrNotKnownFlagsPReg_4_3,storeAddrNotKnownFlagsPReg_4_2,storeAddrNotKnownFlagsPReg_4_1,storeAddrNotKnownFlagsPReg_4_0}; // @[LoadQueue.scala 238:58:@9039.8]
  assign _T_25058 = {lastConflict_4_7,lastConflict_4_6,lastConflict_4_5,lastConflict_4_4,lastConflict_4_3,lastConflict_4_2,lastConflict_4_1,lastConflict_4_0}; // @[LoadQueue.scala 238:96:@9046.8]
  assign _T_25059 = _T_25051 < _T_25058; // @[LoadQueue.scala 238:61:@9047.8]
  assign _T_25060 = canBypass_4 & _T_25059; // @[LoadQueue.scala 237:64:@9048.8]
  assign _GEN_553 = _T_25021 ? _T_25060 : 1'h0; // @[LoadQueue.scala 230:110:@9012.6]
  assign bypassRequest_4 = _T_25013 ? _GEN_553 : 1'h0; // @[LoadQueue.scala 229:71:@9006.4]
  assign _GEN_528 = bypassRequest_4 ? 1'h1 : bypassInitiated_4; // @[LoadQueue.scala 217:34:@8778.6]
  assign _GEN_529 = initBits_4 ? 1'h0 : _GEN_528; // @[LoadQueue.scala 215:23:@8774.4]
  assign _T_25103 = {storeAddrNotKnownFlagsPReg_5_7,storeAddrNotKnownFlagsPReg_5_6,storeAddrNotKnownFlagsPReg_5_5,storeAddrNotKnownFlagsPReg_5_4,storeAddrNotKnownFlagsPReg_5_3,storeAddrNotKnownFlagsPReg_5_2,storeAddrNotKnownFlagsPReg_5_1,storeAddrNotKnownFlagsPReg_5_0}; // @[LoadQueue.scala 238:58:@9089.8]
  assign _T_25110 = {lastConflict_5_7,lastConflict_5_6,lastConflict_5_5,lastConflict_5_4,lastConflict_5_3,lastConflict_5_2,lastConflict_5_1,lastConflict_5_0}; // @[LoadQueue.scala 238:96:@9096.8]
  assign _T_25111 = _T_25103 < _T_25110; // @[LoadQueue.scala 238:61:@9097.8]
  assign _T_25112 = canBypass_5 & _T_25111; // @[LoadQueue.scala 237:64:@9098.8]
  assign _GEN_557 = _T_25073 ? _T_25112 : 1'h0; // @[LoadQueue.scala 230:110:@9062.6]
  assign bypassRequest_5 = _T_25065 ? _GEN_557 : 1'h0; // @[LoadQueue.scala 229:71:@9056.4]
  assign _GEN_530 = bypassRequest_5 ? 1'h1 : bypassInitiated_5; // @[LoadQueue.scala 217:34:@8785.6]
  assign _GEN_531 = initBits_5 ? 1'h0 : _GEN_530; // @[LoadQueue.scala 215:23:@8781.4]
  assign _T_25155 = {storeAddrNotKnownFlagsPReg_6_7,storeAddrNotKnownFlagsPReg_6_6,storeAddrNotKnownFlagsPReg_6_5,storeAddrNotKnownFlagsPReg_6_4,storeAddrNotKnownFlagsPReg_6_3,storeAddrNotKnownFlagsPReg_6_2,storeAddrNotKnownFlagsPReg_6_1,storeAddrNotKnownFlagsPReg_6_0}; // @[LoadQueue.scala 238:58:@9139.8]
  assign _T_25162 = {lastConflict_6_7,lastConflict_6_6,lastConflict_6_5,lastConflict_6_4,lastConflict_6_3,lastConflict_6_2,lastConflict_6_1,lastConflict_6_0}; // @[LoadQueue.scala 238:96:@9146.8]
  assign _T_25163 = _T_25155 < _T_25162; // @[LoadQueue.scala 238:61:@9147.8]
  assign _T_25164 = canBypass_6 & _T_25163; // @[LoadQueue.scala 237:64:@9148.8]
  assign _GEN_561 = _T_25125 ? _T_25164 : 1'h0; // @[LoadQueue.scala 230:110:@9112.6]
  assign bypassRequest_6 = _T_25117 ? _GEN_561 : 1'h0; // @[LoadQueue.scala 229:71:@9106.4]
  assign _GEN_532 = bypassRequest_6 ? 1'h1 : bypassInitiated_6; // @[LoadQueue.scala 217:34:@8792.6]
  assign _GEN_533 = initBits_6 ? 1'h0 : _GEN_532; // @[LoadQueue.scala 215:23:@8788.4]
  assign _T_25207 = {storeAddrNotKnownFlagsPReg_7_7,storeAddrNotKnownFlagsPReg_7_6,storeAddrNotKnownFlagsPReg_7_5,storeAddrNotKnownFlagsPReg_7_4,storeAddrNotKnownFlagsPReg_7_3,storeAddrNotKnownFlagsPReg_7_2,storeAddrNotKnownFlagsPReg_7_1,storeAddrNotKnownFlagsPReg_7_0}; // @[LoadQueue.scala 238:58:@9189.8]
  assign _T_25214 = {lastConflict_7_7,lastConflict_7_6,lastConflict_7_5,lastConflict_7_4,lastConflict_7_3,lastConflict_7_2,lastConflict_7_1,lastConflict_7_0}; // @[LoadQueue.scala 238:96:@9196.8]
  assign _T_25215 = _T_25207 < _T_25214; // @[LoadQueue.scala 238:61:@9197.8]
  assign _T_25216 = canBypass_7 & _T_25215; // @[LoadQueue.scala 237:64:@9198.8]
  assign _GEN_565 = _T_25177 ? _T_25216 : 1'h0; // @[LoadQueue.scala 230:110:@9162.6]
  assign bypassRequest_7 = _T_25169 ? _GEN_565 : 1'h0; // @[LoadQueue.scala 229:71:@9156.4]
  assign _GEN_534 = bypassRequest_7 ? 1'h1 : bypassInitiated_7; // @[LoadQueue.scala 217:34:@8799.6]
  assign _GEN_535 = initBits_7 ? 1'h0 : _GEN_534; // @[LoadQueue.scala 215:23:@8795.4]
  assign _T_25220 = loadRequest_0 | loadRequest_1; // @[LoadQueue.scala 247:28:@9204.4]
  assign _T_25221 = _T_25220 | loadRequest_2; // @[LoadQueue.scala 247:28:@9205.4]
  assign _T_25222 = _T_25221 | loadRequest_3; // @[LoadQueue.scala 247:28:@9206.4]
  assign _T_25223 = _T_25222 | loadRequest_4; // @[LoadQueue.scala 247:28:@9207.4]
  assign _T_25224 = _T_25223 | loadRequest_5; // @[LoadQueue.scala 247:28:@9208.4]
  assign _T_25225 = _T_25224 | loadRequest_6; // @[LoadQueue.scala 247:28:@9209.4]
  assign _T_25226 = _T_25225 | loadRequest_7; // @[LoadQueue.scala 247:28:@9210.4]
  assign _T_25235 = priorityLoadRequest_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@9212.6]
  assign _T_25236 = priorityLoadRequest_5 ? 3'h5 : _T_25235; // @[Mux.scala 31:69:@9213.6]
  assign _T_25237 = priorityLoadRequest_4 ? 3'h4 : _T_25236; // @[Mux.scala 31:69:@9214.6]
  assign _T_25238 = priorityLoadRequest_3 ? 3'h3 : _T_25237; // @[Mux.scala 31:69:@9215.6]
  assign _T_25239 = priorityLoadRequest_2 ? 3'h2 : _T_25238; // @[Mux.scala 31:69:@9216.6]
  assign _T_25240 = priorityLoadRequest_1 ? 3'h1 : _T_25239; // @[Mux.scala 31:69:@9217.6]
  assign _T_25241 = priorityLoadRequest_0 ? 3'h0 : _T_25240; // @[Mux.scala 31:69:@9218.6]
  assign _GEN_569 = 3'h1 == _T_25241 ? addrQ_1 : addrQ_0; // @[LoadQueue.scala 248:24:@9219.6]
  assign _GEN_570 = 3'h2 == _T_25241 ? addrQ_2 : _GEN_569; // @[LoadQueue.scala 248:24:@9219.6]
  assign _GEN_571 = 3'h3 == _T_25241 ? addrQ_3 : _GEN_570; // @[LoadQueue.scala 248:24:@9219.6]
  assign _GEN_572 = 3'h4 == _T_25241 ? addrQ_4 : _GEN_571; // @[LoadQueue.scala 248:24:@9219.6]
  assign _GEN_573 = 3'h5 == _T_25241 ? addrQ_5 : _GEN_572; // @[LoadQueue.scala 248:24:@9219.6]
  assign _GEN_574 = 3'h6 == _T_25241 ? addrQ_6 : _GEN_573; // @[LoadQueue.scala 248:24:@9219.6]
  assign _GEN_575 = 3'h7 == _T_25241 ? addrQ_7 : _GEN_574; // @[LoadQueue.scala 248:24:@9219.6]
  assign _T_25249 = prevPriorityRequest_0 | bypassRequest_0; // @[LoadQueue.scala 261:41:@9230.6]
  assign _GEN_578 = _T_25249 ? 1'h1 : dataKnown_0; // @[LoadQueue.scala 261:62:@9231.6]
  assign _GEN_579 = initBits_0 ? 1'h0 : _GEN_578; // @[LoadQueue.scala 259:25:@9226.4]
  assign _T_25252 = prevPriorityRequest_1 | bypassRequest_1; // @[LoadQueue.scala 261:41:@9238.6]
  assign _GEN_580 = _T_25252 ? 1'h1 : dataKnown_1; // @[LoadQueue.scala 261:62:@9239.6]
  assign _GEN_581 = initBits_1 ? 1'h0 : _GEN_580; // @[LoadQueue.scala 259:25:@9234.4]
  assign _T_25255 = prevPriorityRequest_2 | bypassRequest_2; // @[LoadQueue.scala 261:41:@9246.6]
  assign _GEN_582 = _T_25255 ? 1'h1 : dataKnown_2; // @[LoadQueue.scala 261:62:@9247.6]
  assign _GEN_583 = initBits_2 ? 1'h0 : _GEN_582; // @[LoadQueue.scala 259:25:@9242.4]
  assign _T_25258 = prevPriorityRequest_3 | bypassRequest_3; // @[LoadQueue.scala 261:41:@9254.6]
  assign _GEN_584 = _T_25258 ? 1'h1 : dataKnown_3; // @[LoadQueue.scala 261:62:@9255.6]
  assign _GEN_585 = initBits_3 ? 1'h0 : _GEN_584; // @[LoadQueue.scala 259:25:@9250.4]
  assign _T_25261 = prevPriorityRequest_4 | bypassRequest_4; // @[LoadQueue.scala 261:41:@9262.6]
  assign _GEN_586 = _T_25261 ? 1'h1 : dataKnown_4; // @[LoadQueue.scala 261:62:@9263.6]
  assign _GEN_587 = initBits_4 ? 1'h0 : _GEN_586; // @[LoadQueue.scala 259:25:@9258.4]
  assign _T_25264 = prevPriorityRequest_5 | bypassRequest_5; // @[LoadQueue.scala 261:41:@9270.6]
  assign _GEN_588 = _T_25264 ? 1'h1 : dataKnown_5; // @[LoadQueue.scala 261:62:@9271.6]
  assign _GEN_589 = initBits_5 ? 1'h0 : _GEN_588; // @[LoadQueue.scala 259:25:@9266.4]
  assign _T_25267 = prevPriorityRequest_6 | bypassRequest_6; // @[LoadQueue.scala 261:41:@9278.6]
  assign _GEN_590 = _T_25267 ? 1'h1 : dataKnown_6; // @[LoadQueue.scala 261:62:@9279.6]
  assign _GEN_591 = initBits_6 ? 1'h0 : _GEN_590; // @[LoadQueue.scala 259:25:@9274.4]
  assign _T_25270 = prevPriorityRequest_7 | bypassRequest_7; // @[LoadQueue.scala 261:41:@9286.6]
  assign _GEN_592 = _T_25270 ? 1'h1 : dataKnown_7; // @[LoadQueue.scala 261:62:@9287.6]
  assign _GEN_593 = initBits_7 ? 1'h0 : _GEN_592; // @[LoadQueue.scala 259:25:@9282.4]
  assign _GEN_594 = prevPriorityRequest_0 ? io_loadDataFromMem : dataQ_0; // @[LoadQueue.scala 269:44:@9294.6]
  assign _GEN_595 = bypassRequest_0 ? bypassVal_0 : _GEN_594; // @[LoadQueue.scala 267:32:@9290.4]
  assign _GEN_596 = prevPriorityRequest_1 ? io_loadDataFromMem : dataQ_1; // @[LoadQueue.scala 269:44:@9301.6]
  assign _GEN_597 = bypassRequest_1 ? bypassVal_1 : _GEN_596; // @[LoadQueue.scala 267:32:@9297.4]
  assign _GEN_598 = prevPriorityRequest_2 ? io_loadDataFromMem : dataQ_2; // @[LoadQueue.scala 269:44:@9308.6]
  assign _GEN_599 = bypassRequest_2 ? bypassVal_2 : _GEN_598; // @[LoadQueue.scala 267:32:@9304.4]
  assign _GEN_600 = prevPriorityRequest_3 ? io_loadDataFromMem : dataQ_3; // @[LoadQueue.scala 269:44:@9315.6]
  assign _GEN_601 = bypassRequest_3 ? bypassVal_3 : _GEN_600; // @[LoadQueue.scala 267:32:@9311.4]
  assign _GEN_602 = prevPriorityRequest_4 ? io_loadDataFromMem : dataQ_4; // @[LoadQueue.scala 269:44:@9322.6]
  assign _GEN_603 = bypassRequest_4 ? bypassVal_4 : _GEN_602; // @[LoadQueue.scala 267:32:@9318.4]
  assign _GEN_604 = prevPriorityRequest_5 ? io_loadDataFromMem : dataQ_5; // @[LoadQueue.scala 269:44:@9329.6]
  assign _GEN_605 = bypassRequest_5 ? bypassVal_5 : _GEN_604; // @[LoadQueue.scala 267:32:@9325.4]
  assign _GEN_606 = prevPriorityRequest_6 ? io_loadDataFromMem : dataQ_6; // @[LoadQueue.scala 269:44:@9336.6]
  assign _GEN_607 = bypassRequest_6 ? bypassVal_6 : _GEN_606; // @[LoadQueue.scala 267:32:@9332.4]
  assign _GEN_608 = prevPriorityRequest_7 ? io_loadDataFromMem : dataQ_7; // @[LoadQueue.scala 269:44:@9343.6]
  assign _GEN_609 = bypassRequest_7 ? bypassVal_7 : _GEN_608; // @[LoadQueue.scala 267:32:@9339.4]
  assign entriesPorts_0_0 = portQ_0 == 3'h0; // @[LoadQueue.scala 286:69:@9347.4]
  assign entriesPorts_0_1 = portQ_1 == 3'h0; // @[LoadQueue.scala 286:69:@9349.4]
  assign entriesPorts_0_2 = portQ_2 == 3'h0; // @[LoadQueue.scala 286:69:@9351.4]
  assign entriesPorts_0_3 = portQ_3 == 3'h0; // @[LoadQueue.scala 286:69:@9353.4]
  assign entriesPorts_0_4 = portQ_4 == 3'h0; // @[LoadQueue.scala 286:69:@9355.4]
  assign entriesPorts_0_5 = portQ_5 == 3'h0; // @[LoadQueue.scala 286:69:@9357.4]
  assign entriesPorts_0_6 = portQ_6 == 3'h0; // @[LoadQueue.scala 286:69:@9359.4]
  assign entriesPorts_0_7 = portQ_7 == 3'h0; // @[LoadQueue.scala 286:69:@9361.4]
  assign entriesPorts_1_0 = portQ_0 == 3'h1; // @[LoadQueue.scala 286:69:@9363.4]
  assign entriesPorts_1_1 = portQ_1 == 3'h1; // @[LoadQueue.scala 286:69:@9365.4]
  assign entriesPorts_1_2 = portQ_2 == 3'h1; // @[LoadQueue.scala 286:69:@9367.4]
  assign entriesPorts_1_3 = portQ_3 == 3'h1; // @[LoadQueue.scala 286:69:@9369.4]
  assign entriesPorts_1_4 = portQ_4 == 3'h1; // @[LoadQueue.scala 286:69:@9371.4]
  assign entriesPorts_1_5 = portQ_5 == 3'h1; // @[LoadQueue.scala 286:69:@9373.4]
  assign entriesPorts_1_6 = portQ_6 == 3'h1; // @[LoadQueue.scala 286:69:@9375.4]
  assign entriesPorts_1_7 = portQ_7 == 3'h1; // @[LoadQueue.scala 286:69:@9377.4]
  assign entriesPorts_2_0 = portQ_0 == 3'h2; // @[LoadQueue.scala 286:69:@9379.4]
  assign entriesPorts_2_1 = portQ_1 == 3'h2; // @[LoadQueue.scala 286:69:@9381.4]
  assign entriesPorts_2_2 = portQ_2 == 3'h2; // @[LoadQueue.scala 286:69:@9383.4]
  assign entriesPorts_2_3 = portQ_3 == 3'h2; // @[LoadQueue.scala 286:69:@9385.4]
  assign entriesPorts_2_4 = portQ_4 == 3'h2; // @[LoadQueue.scala 286:69:@9387.4]
  assign entriesPorts_2_5 = portQ_5 == 3'h2; // @[LoadQueue.scala 286:69:@9389.4]
  assign entriesPorts_2_6 = portQ_6 == 3'h2; // @[LoadQueue.scala 286:69:@9391.4]
  assign entriesPorts_2_7 = portQ_7 == 3'h2; // @[LoadQueue.scala 286:69:@9393.4]
  assign entriesPorts_3_0 = portQ_0 == 3'h3; // @[LoadQueue.scala 286:69:@9395.4]
  assign entriesPorts_3_1 = portQ_1 == 3'h3; // @[LoadQueue.scala 286:69:@9397.4]
  assign entriesPorts_3_2 = portQ_2 == 3'h3; // @[LoadQueue.scala 286:69:@9399.4]
  assign entriesPorts_3_3 = portQ_3 == 3'h3; // @[LoadQueue.scala 286:69:@9401.4]
  assign entriesPorts_3_4 = portQ_4 == 3'h3; // @[LoadQueue.scala 286:69:@9403.4]
  assign entriesPorts_3_5 = portQ_5 == 3'h3; // @[LoadQueue.scala 286:69:@9405.4]
  assign entriesPorts_3_6 = portQ_6 == 3'h3; // @[LoadQueue.scala 286:69:@9407.4]
  assign entriesPorts_3_7 = portQ_7 == 3'h3; // @[LoadQueue.scala 286:69:@9409.4]
  assign entriesPorts_4_0 = portQ_0 == 3'h4; // @[LoadQueue.scala 286:69:@9411.4]
  assign entriesPorts_4_1 = portQ_1 == 3'h4; // @[LoadQueue.scala 286:69:@9413.4]
  assign entriesPorts_4_2 = portQ_2 == 3'h4; // @[LoadQueue.scala 286:69:@9415.4]
  assign entriesPorts_4_3 = portQ_3 == 3'h4; // @[LoadQueue.scala 286:69:@9417.4]
  assign entriesPorts_4_4 = portQ_4 == 3'h4; // @[LoadQueue.scala 286:69:@9419.4]
  assign entriesPorts_4_5 = portQ_5 == 3'h4; // @[LoadQueue.scala 286:69:@9421.4]
  assign entriesPorts_4_6 = portQ_6 == 3'h4; // @[LoadQueue.scala 286:69:@9423.4]
  assign entriesPorts_4_7 = portQ_7 == 3'h4; // @[LoadQueue.scala 286:69:@9425.4]
  assign _T_26091 = addrKnown_0 == 1'h0; // @[LoadQueue.scala 298:86:@9429.4]
  assign _T_26092 = entriesPorts_0_0 & _T_26091; // @[LoadQueue.scala 298:83:@9430.4]
  assign _T_26094 = addrKnown_1 == 1'h0; // @[LoadQueue.scala 298:86:@9431.4]
  assign _T_26095 = entriesPorts_0_1 & _T_26094; // @[LoadQueue.scala 298:83:@9432.4]
  assign _T_26097 = addrKnown_2 == 1'h0; // @[LoadQueue.scala 298:86:@9433.4]
  assign _T_26098 = entriesPorts_0_2 & _T_26097; // @[LoadQueue.scala 298:83:@9434.4]
  assign _T_26100 = addrKnown_3 == 1'h0; // @[LoadQueue.scala 298:86:@9435.4]
  assign _T_26101 = entriesPorts_0_3 & _T_26100; // @[LoadQueue.scala 298:83:@9436.4]
  assign _T_26103 = addrKnown_4 == 1'h0; // @[LoadQueue.scala 298:86:@9437.4]
  assign _T_26104 = entriesPorts_0_4 & _T_26103; // @[LoadQueue.scala 298:83:@9438.4]
  assign _T_26106 = addrKnown_5 == 1'h0; // @[LoadQueue.scala 298:86:@9439.4]
  assign _T_26107 = entriesPorts_0_5 & _T_26106; // @[LoadQueue.scala 298:83:@9440.4]
  assign _T_26109 = addrKnown_6 == 1'h0; // @[LoadQueue.scala 298:86:@9441.4]
  assign _T_26110 = entriesPorts_0_6 & _T_26109; // @[LoadQueue.scala 298:83:@9442.4]
  assign _T_26112 = addrKnown_7 == 1'h0; // @[LoadQueue.scala 298:86:@9443.4]
  assign _T_26113 = entriesPorts_0_7 & _T_26112; // @[LoadQueue.scala 298:83:@9444.4]
  assign _T_26164 = _T_26113 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9474.4]
  assign _T_26165 = _T_26110 ? 8'h40 : _T_26164; // @[Mux.scala 31:69:@9475.4]
  assign _T_26166 = _T_26107 ? 8'h20 : _T_26165; // @[Mux.scala 31:69:@9476.4]
  assign _T_26167 = _T_26104 ? 8'h10 : _T_26166; // @[Mux.scala 31:69:@9477.4]
  assign _T_26168 = _T_26101 ? 8'h8 : _T_26167; // @[Mux.scala 31:69:@9478.4]
  assign _T_26169 = _T_26098 ? 8'h4 : _T_26168; // @[Mux.scala 31:69:@9479.4]
  assign _T_26170 = _T_26095 ? 8'h2 : _T_26169; // @[Mux.scala 31:69:@9480.4]
  assign _T_26171 = _T_26092 ? 8'h1 : _T_26170; // @[Mux.scala 31:69:@9481.4]
  assign _T_26172 = _T_26171[0]; // @[OneHot.scala 66:30:@9482.4]
  assign _T_26173 = _T_26171[1]; // @[OneHot.scala 66:30:@9483.4]
  assign _T_26174 = _T_26171[2]; // @[OneHot.scala 66:30:@9484.4]
  assign _T_26175 = _T_26171[3]; // @[OneHot.scala 66:30:@9485.4]
  assign _T_26176 = _T_26171[4]; // @[OneHot.scala 66:30:@9486.4]
  assign _T_26177 = _T_26171[5]; // @[OneHot.scala 66:30:@9487.4]
  assign _T_26178 = _T_26171[6]; // @[OneHot.scala 66:30:@9488.4]
  assign _T_26179 = _T_26171[7]; // @[OneHot.scala 66:30:@9489.4]
  assign _T_26204 = _T_26092 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9499.4]
  assign _T_26205 = _T_26113 ? 8'h40 : _T_26204; // @[Mux.scala 31:69:@9500.4]
  assign _T_26206 = _T_26110 ? 8'h20 : _T_26205; // @[Mux.scala 31:69:@9501.4]
  assign _T_26207 = _T_26107 ? 8'h10 : _T_26206; // @[Mux.scala 31:69:@9502.4]
  assign _T_26208 = _T_26104 ? 8'h8 : _T_26207; // @[Mux.scala 31:69:@9503.4]
  assign _T_26209 = _T_26101 ? 8'h4 : _T_26208; // @[Mux.scala 31:69:@9504.4]
  assign _T_26210 = _T_26098 ? 8'h2 : _T_26209; // @[Mux.scala 31:69:@9505.4]
  assign _T_26211 = _T_26095 ? 8'h1 : _T_26210; // @[Mux.scala 31:69:@9506.4]
  assign _T_26212 = _T_26211[0]; // @[OneHot.scala 66:30:@9507.4]
  assign _T_26213 = _T_26211[1]; // @[OneHot.scala 66:30:@9508.4]
  assign _T_26214 = _T_26211[2]; // @[OneHot.scala 66:30:@9509.4]
  assign _T_26215 = _T_26211[3]; // @[OneHot.scala 66:30:@9510.4]
  assign _T_26216 = _T_26211[4]; // @[OneHot.scala 66:30:@9511.4]
  assign _T_26217 = _T_26211[5]; // @[OneHot.scala 66:30:@9512.4]
  assign _T_26218 = _T_26211[6]; // @[OneHot.scala 66:30:@9513.4]
  assign _T_26219 = _T_26211[7]; // @[OneHot.scala 66:30:@9514.4]
  assign _T_26244 = _T_26095 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9524.4]
  assign _T_26245 = _T_26092 ? 8'h40 : _T_26244; // @[Mux.scala 31:69:@9525.4]
  assign _T_26246 = _T_26113 ? 8'h20 : _T_26245; // @[Mux.scala 31:69:@9526.4]
  assign _T_26247 = _T_26110 ? 8'h10 : _T_26246; // @[Mux.scala 31:69:@9527.4]
  assign _T_26248 = _T_26107 ? 8'h8 : _T_26247; // @[Mux.scala 31:69:@9528.4]
  assign _T_26249 = _T_26104 ? 8'h4 : _T_26248; // @[Mux.scala 31:69:@9529.4]
  assign _T_26250 = _T_26101 ? 8'h2 : _T_26249; // @[Mux.scala 31:69:@9530.4]
  assign _T_26251 = _T_26098 ? 8'h1 : _T_26250; // @[Mux.scala 31:69:@9531.4]
  assign _T_26252 = _T_26251[0]; // @[OneHot.scala 66:30:@9532.4]
  assign _T_26253 = _T_26251[1]; // @[OneHot.scala 66:30:@9533.4]
  assign _T_26254 = _T_26251[2]; // @[OneHot.scala 66:30:@9534.4]
  assign _T_26255 = _T_26251[3]; // @[OneHot.scala 66:30:@9535.4]
  assign _T_26256 = _T_26251[4]; // @[OneHot.scala 66:30:@9536.4]
  assign _T_26257 = _T_26251[5]; // @[OneHot.scala 66:30:@9537.4]
  assign _T_26258 = _T_26251[6]; // @[OneHot.scala 66:30:@9538.4]
  assign _T_26259 = _T_26251[7]; // @[OneHot.scala 66:30:@9539.4]
  assign _T_26284 = _T_26098 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9549.4]
  assign _T_26285 = _T_26095 ? 8'h40 : _T_26284; // @[Mux.scala 31:69:@9550.4]
  assign _T_26286 = _T_26092 ? 8'h20 : _T_26285; // @[Mux.scala 31:69:@9551.4]
  assign _T_26287 = _T_26113 ? 8'h10 : _T_26286; // @[Mux.scala 31:69:@9552.4]
  assign _T_26288 = _T_26110 ? 8'h8 : _T_26287; // @[Mux.scala 31:69:@9553.4]
  assign _T_26289 = _T_26107 ? 8'h4 : _T_26288; // @[Mux.scala 31:69:@9554.4]
  assign _T_26290 = _T_26104 ? 8'h2 : _T_26289; // @[Mux.scala 31:69:@9555.4]
  assign _T_26291 = _T_26101 ? 8'h1 : _T_26290; // @[Mux.scala 31:69:@9556.4]
  assign _T_26292 = _T_26291[0]; // @[OneHot.scala 66:30:@9557.4]
  assign _T_26293 = _T_26291[1]; // @[OneHot.scala 66:30:@9558.4]
  assign _T_26294 = _T_26291[2]; // @[OneHot.scala 66:30:@9559.4]
  assign _T_26295 = _T_26291[3]; // @[OneHot.scala 66:30:@9560.4]
  assign _T_26296 = _T_26291[4]; // @[OneHot.scala 66:30:@9561.4]
  assign _T_26297 = _T_26291[5]; // @[OneHot.scala 66:30:@9562.4]
  assign _T_26298 = _T_26291[6]; // @[OneHot.scala 66:30:@9563.4]
  assign _T_26299 = _T_26291[7]; // @[OneHot.scala 66:30:@9564.4]
  assign _T_26324 = _T_26101 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9574.4]
  assign _T_26325 = _T_26098 ? 8'h40 : _T_26324; // @[Mux.scala 31:69:@9575.4]
  assign _T_26326 = _T_26095 ? 8'h20 : _T_26325; // @[Mux.scala 31:69:@9576.4]
  assign _T_26327 = _T_26092 ? 8'h10 : _T_26326; // @[Mux.scala 31:69:@9577.4]
  assign _T_26328 = _T_26113 ? 8'h8 : _T_26327; // @[Mux.scala 31:69:@9578.4]
  assign _T_26329 = _T_26110 ? 8'h4 : _T_26328; // @[Mux.scala 31:69:@9579.4]
  assign _T_26330 = _T_26107 ? 8'h2 : _T_26329; // @[Mux.scala 31:69:@9580.4]
  assign _T_26331 = _T_26104 ? 8'h1 : _T_26330; // @[Mux.scala 31:69:@9581.4]
  assign _T_26332 = _T_26331[0]; // @[OneHot.scala 66:30:@9582.4]
  assign _T_26333 = _T_26331[1]; // @[OneHot.scala 66:30:@9583.4]
  assign _T_26334 = _T_26331[2]; // @[OneHot.scala 66:30:@9584.4]
  assign _T_26335 = _T_26331[3]; // @[OneHot.scala 66:30:@9585.4]
  assign _T_26336 = _T_26331[4]; // @[OneHot.scala 66:30:@9586.4]
  assign _T_26337 = _T_26331[5]; // @[OneHot.scala 66:30:@9587.4]
  assign _T_26338 = _T_26331[6]; // @[OneHot.scala 66:30:@9588.4]
  assign _T_26339 = _T_26331[7]; // @[OneHot.scala 66:30:@9589.4]
  assign _T_26364 = _T_26104 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9599.4]
  assign _T_26365 = _T_26101 ? 8'h40 : _T_26364; // @[Mux.scala 31:69:@9600.4]
  assign _T_26366 = _T_26098 ? 8'h20 : _T_26365; // @[Mux.scala 31:69:@9601.4]
  assign _T_26367 = _T_26095 ? 8'h10 : _T_26366; // @[Mux.scala 31:69:@9602.4]
  assign _T_26368 = _T_26092 ? 8'h8 : _T_26367; // @[Mux.scala 31:69:@9603.4]
  assign _T_26369 = _T_26113 ? 8'h4 : _T_26368; // @[Mux.scala 31:69:@9604.4]
  assign _T_26370 = _T_26110 ? 8'h2 : _T_26369; // @[Mux.scala 31:69:@9605.4]
  assign _T_26371 = _T_26107 ? 8'h1 : _T_26370; // @[Mux.scala 31:69:@9606.4]
  assign _T_26372 = _T_26371[0]; // @[OneHot.scala 66:30:@9607.4]
  assign _T_26373 = _T_26371[1]; // @[OneHot.scala 66:30:@9608.4]
  assign _T_26374 = _T_26371[2]; // @[OneHot.scala 66:30:@9609.4]
  assign _T_26375 = _T_26371[3]; // @[OneHot.scala 66:30:@9610.4]
  assign _T_26376 = _T_26371[4]; // @[OneHot.scala 66:30:@9611.4]
  assign _T_26377 = _T_26371[5]; // @[OneHot.scala 66:30:@9612.4]
  assign _T_26378 = _T_26371[6]; // @[OneHot.scala 66:30:@9613.4]
  assign _T_26379 = _T_26371[7]; // @[OneHot.scala 66:30:@9614.4]
  assign _T_26404 = _T_26107 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9624.4]
  assign _T_26405 = _T_26104 ? 8'h40 : _T_26404; // @[Mux.scala 31:69:@9625.4]
  assign _T_26406 = _T_26101 ? 8'h20 : _T_26405; // @[Mux.scala 31:69:@9626.4]
  assign _T_26407 = _T_26098 ? 8'h10 : _T_26406; // @[Mux.scala 31:69:@9627.4]
  assign _T_26408 = _T_26095 ? 8'h8 : _T_26407; // @[Mux.scala 31:69:@9628.4]
  assign _T_26409 = _T_26092 ? 8'h4 : _T_26408; // @[Mux.scala 31:69:@9629.4]
  assign _T_26410 = _T_26113 ? 8'h2 : _T_26409; // @[Mux.scala 31:69:@9630.4]
  assign _T_26411 = _T_26110 ? 8'h1 : _T_26410; // @[Mux.scala 31:69:@9631.4]
  assign _T_26412 = _T_26411[0]; // @[OneHot.scala 66:30:@9632.4]
  assign _T_26413 = _T_26411[1]; // @[OneHot.scala 66:30:@9633.4]
  assign _T_26414 = _T_26411[2]; // @[OneHot.scala 66:30:@9634.4]
  assign _T_26415 = _T_26411[3]; // @[OneHot.scala 66:30:@9635.4]
  assign _T_26416 = _T_26411[4]; // @[OneHot.scala 66:30:@9636.4]
  assign _T_26417 = _T_26411[5]; // @[OneHot.scala 66:30:@9637.4]
  assign _T_26418 = _T_26411[6]; // @[OneHot.scala 66:30:@9638.4]
  assign _T_26419 = _T_26411[7]; // @[OneHot.scala 66:30:@9639.4]
  assign _T_26444 = _T_26110 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9649.4]
  assign _T_26445 = _T_26107 ? 8'h40 : _T_26444; // @[Mux.scala 31:69:@9650.4]
  assign _T_26446 = _T_26104 ? 8'h20 : _T_26445; // @[Mux.scala 31:69:@9651.4]
  assign _T_26447 = _T_26101 ? 8'h10 : _T_26446; // @[Mux.scala 31:69:@9652.4]
  assign _T_26448 = _T_26098 ? 8'h8 : _T_26447; // @[Mux.scala 31:69:@9653.4]
  assign _T_26449 = _T_26095 ? 8'h4 : _T_26448; // @[Mux.scala 31:69:@9654.4]
  assign _T_26450 = _T_26092 ? 8'h2 : _T_26449; // @[Mux.scala 31:69:@9655.4]
  assign _T_26451 = _T_26113 ? 8'h1 : _T_26450; // @[Mux.scala 31:69:@9656.4]
  assign _T_26452 = _T_26451[0]; // @[OneHot.scala 66:30:@9657.4]
  assign _T_26453 = _T_26451[1]; // @[OneHot.scala 66:30:@9658.4]
  assign _T_26454 = _T_26451[2]; // @[OneHot.scala 66:30:@9659.4]
  assign _T_26455 = _T_26451[3]; // @[OneHot.scala 66:30:@9660.4]
  assign _T_26456 = _T_26451[4]; // @[OneHot.scala 66:30:@9661.4]
  assign _T_26457 = _T_26451[5]; // @[OneHot.scala 66:30:@9662.4]
  assign _T_26458 = _T_26451[6]; // @[OneHot.scala 66:30:@9663.4]
  assign _T_26459 = _T_26451[7]; // @[OneHot.scala 66:30:@9664.4]
  assign _T_26500 = {_T_26179,_T_26178,_T_26177,_T_26176,_T_26175,_T_26174,_T_26173,_T_26172}; // @[Mux.scala 19:72:@9680.4]
  assign _T_26502 = _T_24176 ? _T_26500 : 8'h0; // @[Mux.scala 19:72:@9681.4]
  assign _T_26509 = {_T_26218,_T_26217,_T_26216,_T_26215,_T_26214,_T_26213,_T_26212,_T_26219}; // @[Mux.scala 19:72:@9688.4]
  assign _T_26511 = _T_24177 ? _T_26509 : 8'h0; // @[Mux.scala 19:72:@9689.4]
  assign _T_26518 = {_T_26257,_T_26256,_T_26255,_T_26254,_T_26253,_T_26252,_T_26259,_T_26258}; // @[Mux.scala 19:72:@9696.4]
  assign _T_26520 = _T_24178 ? _T_26518 : 8'h0; // @[Mux.scala 19:72:@9697.4]
  assign _T_26527 = {_T_26296,_T_26295,_T_26294,_T_26293,_T_26292,_T_26299,_T_26298,_T_26297}; // @[Mux.scala 19:72:@9704.4]
  assign _T_26529 = _T_24179 ? _T_26527 : 8'h0; // @[Mux.scala 19:72:@9705.4]
  assign _T_26536 = {_T_26335,_T_26334,_T_26333,_T_26332,_T_26339,_T_26338,_T_26337,_T_26336}; // @[Mux.scala 19:72:@9712.4]
  assign _T_26538 = _T_24180 ? _T_26536 : 8'h0; // @[Mux.scala 19:72:@9713.4]
  assign _T_26545 = {_T_26374,_T_26373,_T_26372,_T_26379,_T_26378,_T_26377,_T_26376,_T_26375}; // @[Mux.scala 19:72:@9720.4]
  assign _T_26547 = _T_24181 ? _T_26545 : 8'h0; // @[Mux.scala 19:72:@9721.4]
  assign _T_26554 = {_T_26413,_T_26412,_T_26419,_T_26418,_T_26417,_T_26416,_T_26415,_T_26414}; // @[Mux.scala 19:72:@9728.4]
  assign _T_26556 = _T_24182 ? _T_26554 : 8'h0; // @[Mux.scala 19:72:@9729.4]
  assign _T_26563 = {_T_26452,_T_26459,_T_26458,_T_26457,_T_26456,_T_26455,_T_26454,_T_26453}; // @[Mux.scala 19:72:@9736.4]
  assign _T_26565 = _T_24183 ? _T_26563 : 8'h0; // @[Mux.scala 19:72:@9737.4]
  assign _T_26566 = _T_26502 | _T_26511; // @[Mux.scala 19:72:@9738.4]
  assign _T_26567 = _T_26566 | _T_26520; // @[Mux.scala 19:72:@9739.4]
  assign _T_26568 = _T_26567 | _T_26529; // @[Mux.scala 19:72:@9740.4]
  assign _T_26569 = _T_26568 | _T_26538; // @[Mux.scala 19:72:@9741.4]
  assign _T_26570 = _T_26569 | _T_26547; // @[Mux.scala 19:72:@9742.4]
  assign _T_26571 = _T_26570 | _T_26556; // @[Mux.scala 19:72:@9743.4]
  assign _T_26572 = _T_26571 | _T_26565; // @[Mux.scala 19:72:@9744.4]
  assign inputPriorityPorts_0_0 = _T_26572[0]; // @[Mux.scala 19:72:@9748.4]
  assign inputPriorityPorts_0_1 = _T_26572[1]; // @[Mux.scala 19:72:@9750.4]
  assign inputPriorityPorts_0_2 = _T_26572[2]; // @[Mux.scala 19:72:@9752.4]
  assign inputPriorityPorts_0_3 = _T_26572[3]; // @[Mux.scala 19:72:@9754.4]
  assign inputPriorityPorts_0_4 = _T_26572[4]; // @[Mux.scala 19:72:@9756.4]
  assign inputPriorityPorts_0_5 = _T_26572[5]; // @[Mux.scala 19:72:@9758.4]
  assign inputPriorityPorts_0_6 = _T_26572[6]; // @[Mux.scala 19:72:@9760.4]
  assign inputPriorityPorts_0_7 = _T_26572[7]; // @[Mux.scala 19:72:@9762.4]
  assign _T_26686 = entriesPorts_0_7 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9792.4]
  assign _T_26687 = entriesPorts_0_6 ? 8'h40 : _T_26686; // @[Mux.scala 31:69:@9793.4]
  assign _T_26688 = entriesPorts_0_5 ? 8'h20 : _T_26687; // @[Mux.scala 31:69:@9794.4]
  assign _T_26689 = entriesPorts_0_4 ? 8'h10 : _T_26688; // @[Mux.scala 31:69:@9795.4]
  assign _T_26690 = entriesPorts_0_3 ? 8'h8 : _T_26689; // @[Mux.scala 31:69:@9796.4]
  assign _T_26691 = entriesPorts_0_2 ? 8'h4 : _T_26690; // @[Mux.scala 31:69:@9797.4]
  assign _T_26692 = entriesPorts_0_1 ? 8'h2 : _T_26691; // @[Mux.scala 31:69:@9798.4]
  assign _T_26693 = entriesPorts_0_0 ? 8'h1 : _T_26692; // @[Mux.scala 31:69:@9799.4]
  assign _T_26694 = _T_26693[0]; // @[OneHot.scala 66:30:@9800.4]
  assign _T_26695 = _T_26693[1]; // @[OneHot.scala 66:30:@9801.4]
  assign _T_26696 = _T_26693[2]; // @[OneHot.scala 66:30:@9802.4]
  assign _T_26697 = _T_26693[3]; // @[OneHot.scala 66:30:@9803.4]
  assign _T_26698 = _T_26693[4]; // @[OneHot.scala 66:30:@9804.4]
  assign _T_26699 = _T_26693[5]; // @[OneHot.scala 66:30:@9805.4]
  assign _T_26700 = _T_26693[6]; // @[OneHot.scala 66:30:@9806.4]
  assign _T_26701 = _T_26693[7]; // @[OneHot.scala 66:30:@9807.4]
  assign _T_26726 = entriesPorts_0_0 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9817.4]
  assign _T_26727 = entriesPorts_0_7 ? 8'h40 : _T_26726; // @[Mux.scala 31:69:@9818.4]
  assign _T_26728 = entriesPorts_0_6 ? 8'h20 : _T_26727; // @[Mux.scala 31:69:@9819.4]
  assign _T_26729 = entriesPorts_0_5 ? 8'h10 : _T_26728; // @[Mux.scala 31:69:@9820.4]
  assign _T_26730 = entriesPorts_0_4 ? 8'h8 : _T_26729; // @[Mux.scala 31:69:@9821.4]
  assign _T_26731 = entriesPorts_0_3 ? 8'h4 : _T_26730; // @[Mux.scala 31:69:@9822.4]
  assign _T_26732 = entriesPorts_0_2 ? 8'h2 : _T_26731; // @[Mux.scala 31:69:@9823.4]
  assign _T_26733 = entriesPorts_0_1 ? 8'h1 : _T_26732; // @[Mux.scala 31:69:@9824.4]
  assign _T_26734 = _T_26733[0]; // @[OneHot.scala 66:30:@9825.4]
  assign _T_26735 = _T_26733[1]; // @[OneHot.scala 66:30:@9826.4]
  assign _T_26736 = _T_26733[2]; // @[OneHot.scala 66:30:@9827.4]
  assign _T_26737 = _T_26733[3]; // @[OneHot.scala 66:30:@9828.4]
  assign _T_26738 = _T_26733[4]; // @[OneHot.scala 66:30:@9829.4]
  assign _T_26739 = _T_26733[5]; // @[OneHot.scala 66:30:@9830.4]
  assign _T_26740 = _T_26733[6]; // @[OneHot.scala 66:30:@9831.4]
  assign _T_26741 = _T_26733[7]; // @[OneHot.scala 66:30:@9832.4]
  assign _T_26766 = entriesPorts_0_1 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9842.4]
  assign _T_26767 = entriesPorts_0_0 ? 8'h40 : _T_26766; // @[Mux.scala 31:69:@9843.4]
  assign _T_26768 = entriesPorts_0_7 ? 8'h20 : _T_26767; // @[Mux.scala 31:69:@9844.4]
  assign _T_26769 = entriesPorts_0_6 ? 8'h10 : _T_26768; // @[Mux.scala 31:69:@9845.4]
  assign _T_26770 = entriesPorts_0_5 ? 8'h8 : _T_26769; // @[Mux.scala 31:69:@9846.4]
  assign _T_26771 = entriesPorts_0_4 ? 8'h4 : _T_26770; // @[Mux.scala 31:69:@9847.4]
  assign _T_26772 = entriesPorts_0_3 ? 8'h2 : _T_26771; // @[Mux.scala 31:69:@9848.4]
  assign _T_26773 = entriesPorts_0_2 ? 8'h1 : _T_26772; // @[Mux.scala 31:69:@9849.4]
  assign _T_26774 = _T_26773[0]; // @[OneHot.scala 66:30:@9850.4]
  assign _T_26775 = _T_26773[1]; // @[OneHot.scala 66:30:@9851.4]
  assign _T_26776 = _T_26773[2]; // @[OneHot.scala 66:30:@9852.4]
  assign _T_26777 = _T_26773[3]; // @[OneHot.scala 66:30:@9853.4]
  assign _T_26778 = _T_26773[4]; // @[OneHot.scala 66:30:@9854.4]
  assign _T_26779 = _T_26773[5]; // @[OneHot.scala 66:30:@9855.4]
  assign _T_26780 = _T_26773[6]; // @[OneHot.scala 66:30:@9856.4]
  assign _T_26781 = _T_26773[7]; // @[OneHot.scala 66:30:@9857.4]
  assign _T_26806 = entriesPorts_0_2 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9867.4]
  assign _T_26807 = entriesPorts_0_1 ? 8'h40 : _T_26806; // @[Mux.scala 31:69:@9868.4]
  assign _T_26808 = entriesPorts_0_0 ? 8'h20 : _T_26807; // @[Mux.scala 31:69:@9869.4]
  assign _T_26809 = entriesPorts_0_7 ? 8'h10 : _T_26808; // @[Mux.scala 31:69:@9870.4]
  assign _T_26810 = entriesPorts_0_6 ? 8'h8 : _T_26809; // @[Mux.scala 31:69:@9871.4]
  assign _T_26811 = entriesPorts_0_5 ? 8'h4 : _T_26810; // @[Mux.scala 31:69:@9872.4]
  assign _T_26812 = entriesPorts_0_4 ? 8'h2 : _T_26811; // @[Mux.scala 31:69:@9873.4]
  assign _T_26813 = entriesPorts_0_3 ? 8'h1 : _T_26812; // @[Mux.scala 31:69:@9874.4]
  assign _T_26814 = _T_26813[0]; // @[OneHot.scala 66:30:@9875.4]
  assign _T_26815 = _T_26813[1]; // @[OneHot.scala 66:30:@9876.4]
  assign _T_26816 = _T_26813[2]; // @[OneHot.scala 66:30:@9877.4]
  assign _T_26817 = _T_26813[3]; // @[OneHot.scala 66:30:@9878.4]
  assign _T_26818 = _T_26813[4]; // @[OneHot.scala 66:30:@9879.4]
  assign _T_26819 = _T_26813[5]; // @[OneHot.scala 66:30:@9880.4]
  assign _T_26820 = _T_26813[6]; // @[OneHot.scala 66:30:@9881.4]
  assign _T_26821 = _T_26813[7]; // @[OneHot.scala 66:30:@9882.4]
  assign _T_26846 = entriesPorts_0_3 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9892.4]
  assign _T_26847 = entriesPorts_0_2 ? 8'h40 : _T_26846; // @[Mux.scala 31:69:@9893.4]
  assign _T_26848 = entriesPorts_0_1 ? 8'h20 : _T_26847; // @[Mux.scala 31:69:@9894.4]
  assign _T_26849 = entriesPorts_0_0 ? 8'h10 : _T_26848; // @[Mux.scala 31:69:@9895.4]
  assign _T_26850 = entriesPorts_0_7 ? 8'h8 : _T_26849; // @[Mux.scala 31:69:@9896.4]
  assign _T_26851 = entriesPorts_0_6 ? 8'h4 : _T_26850; // @[Mux.scala 31:69:@9897.4]
  assign _T_26852 = entriesPorts_0_5 ? 8'h2 : _T_26851; // @[Mux.scala 31:69:@9898.4]
  assign _T_26853 = entriesPorts_0_4 ? 8'h1 : _T_26852; // @[Mux.scala 31:69:@9899.4]
  assign _T_26854 = _T_26853[0]; // @[OneHot.scala 66:30:@9900.4]
  assign _T_26855 = _T_26853[1]; // @[OneHot.scala 66:30:@9901.4]
  assign _T_26856 = _T_26853[2]; // @[OneHot.scala 66:30:@9902.4]
  assign _T_26857 = _T_26853[3]; // @[OneHot.scala 66:30:@9903.4]
  assign _T_26858 = _T_26853[4]; // @[OneHot.scala 66:30:@9904.4]
  assign _T_26859 = _T_26853[5]; // @[OneHot.scala 66:30:@9905.4]
  assign _T_26860 = _T_26853[6]; // @[OneHot.scala 66:30:@9906.4]
  assign _T_26861 = _T_26853[7]; // @[OneHot.scala 66:30:@9907.4]
  assign _T_26886 = entriesPorts_0_4 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9917.4]
  assign _T_26887 = entriesPorts_0_3 ? 8'h40 : _T_26886; // @[Mux.scala 31:69:@9918.4]
  assign _T_26888 = entriesPorts_0_2 ? 8'h20 : _T_26887; // @[Mux.scala 31:69:@9919.4]
  assign _T_26889 = entriesPorts_0_1 ? 8'h10 : _T_26888; // @[Mux.scala 31:69:@9920.4]
  assign _T_26890 = entriesPorts_0_0 ? 8'h8 : _T_26889; // @[Mux.scala 31:69:@9921.4]
  assign _T_26891 = entriesPorts_0_7 ? 8'h4 : _T_26890; // @[Mux.scala 31:69:@9922.4]
  assign _T_26892 = entriesPorts_0_6 ? 8'h2 : _T_26891; // @[Mux.scala 31:69:@9923.4]
  assign _T_26893 = entriesPorts_0_5 ? 8'h1 : _T_26892; // @[Mux.scala 31:69:@9924.4]
  assign _T_26894 = _T_26893[0]; // @[OneHot.scala 66:30:@9925.4]
  assign _T_26895 = _T_26893[1]; // @[OneHot.scala 66:30:@9926.4]
  assign _T_26896 = _T_26893[2]; // @[OneHot.scala 66:30:@9927.4]
  assign _T_26897 = _T_26893[3]; // @[OneHot.scala 66:30:@9928.4]
  assign _T_26898 = _T_26893[4]; // @[OneHot.scala 66:30:@9929.4]
  assign _T_26899 = _T_26893[5]; // @[OneHot.scala 66:30:@9930.4]
  assign _T_26900 = _T_26893[6]; // @[OneHot.scala 66:30:@9931.4]
  assign _T_26901 = _T_26893[7]; // @[OneHot.scala 66:30:@9932.4]
  assign _T_26926 = entriesPorts_0_5 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9942.4]
  assign _T_26927 = entriesPorts_0_4 ? 8'h40 : _T_26926; // @[Mux.scala 31:69:@9943.4]
  assign _T_26928 = entriesPorts_0_3 ? 8'h20 : _T_26927; // @[Mux.scala 31:69:@9944.4]
  assign _T_26929 = entriesPorts_0_2 ? 8'h10 : _T_26928; // @[Mux.scala 31:69:@9945.4]
  assign _T_26930 = entriesPorts_0_1 ? 8'h8 : _T_26929; // @[Mux.scala 31:69:@9946.4]
  assign _T_26931 = entriesPorts_0_0 ? 8'h4 : _T_26930; // @[Mux.scala 31:69:@9947.4]
  assign _T_26932 = entriesPorts_0_7 ? 8'h2 : _T_26931; // @[Mux.scala 31:69:@9948.4]
  assign _T_26933 = entriesPorts_0_6 ? 8'h1 : _T_26932; // @[Mux.scala 31:69:@9949.4]
  assign _T_26934 = _T_26933[0]; // @[OneHot.scala 66:30:@9950.4]
  assign _T_26935 = _T_26933[1]; // @[OneHot.scala 66:30:@9951.4]
  assign _T_26936 = _T_26933[2]; // @[OneHot.scala 66:30:@9952.4]
  assign _T_26937 = _T_26933[3]; // @[OneHot.scala 66:30:@9953.4]
  assign _T_26938 = _T_26933[4]; // @[OneHot.scala 66:30:@9954.4]
  assign _T_26939 = _T_26933[5]; // @[OneHot.scala 66:30:@9955.4]
  assign _T_26940 = _T_26933[6]; // @[OneHot.scala 66:30:@9956.4]
  assign _T_26941 = _T_26933[7]; // @[OneHot.scala 66:30:@9957.4]
  assign _T_26966 = entriesPorts_0_6 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9967.4]
  assign _T_26967 = entriesPorts_0_5 ? 8'h40 : _T_26966; // @[Mux.scala 31:69:@9968.4]
  assign _T_26968 = entriesPorts_0_4 ? 8'h20 : _T_26967; // @[Mux.scala 31:69:@9969.4]
  assign _T_26969 = entriesPorts_0_3 ? 8'h10 : _T_26968; // @[Mux.scala 31:69:@9970.4]
  assign _T_26970 = entriesPorts_0_2 ? 8'h8 : _T_26969; // @[Mux.scala 31:69:@9971.4]
  assign _T_26971 = entriesPorts_0_1 ? 8'h4 : _T_26970; // @[Mux.scala 31:69:@9972.4]
  assign _T_26972 = entriesPorts_0_0 ? 8'h2 : _T_26971; // @[Mux.scala 31:69:@9973.4]
  assign _T_26973 = entriesPorts_0_7 ? 8'h1 : _T_26972; // @[Mux.scala 31:69:@9974.4]
  assign _T_26974 = _T_26973[0]; // @[OneHot.scala 66:30:@9975.4]
  assign _T_26975 = _T_26973[1]; // @[OneHot.scala 66:30:@9976.4]
  assign _T_26976 = _T_26973[2]; // @[OneHot.scala 66:30:@9977.4]
  assign _T_26977 = _T_26973[3]; // @[OneHot.scala 66:30:@9978.4]
  assign _T_26978 = _T_26973[4]; // @[OneHot.scala 66:30:@9979.4]
  assign _T_26979 = _T_26973[5]; // @[OneHot.scala 66:30:@9980.4]
  assign _T_26980 = _T_26973[6]; // @[OneHot.scala 66:30:@9981.4]
  assign _T_26981 = _T_26973[7]; // @[OneHot.scala 66:30:@9982.4]
  assign _T_27022 = {_T_26701,_T_26700,_T_26699,_T_26698,_T_26697,_T_26696,_T_26695,_T_26694}; // @[Mux.scala 19:72:@9998.4]
  assign _T_27024 = _T_24176 ? _T_27022 : 8'h0; // @[Mux.scala 19:72:@9999.4]
  assign _T_27031 = {_T_26740,_T_26739,_T_26738,_T_26737,_T_26736,_T_26735,_T_26734,_T_26741}; // @[Mux.scala 19:72:@10006.4]
  assign _T_27033 = _T_24177 ? _T_27031 : 8'h0; // @[Mux.scala 19:72:@10007.4]
  assign _T_27040 = {_T_26779,_T_26778,_T_26777,_T_26776,_T_26775,_T_26774,_T_26781,_T_26780}; // @[Mux.scala 19:72:@10014.4]
  assign _T_27042 = _T_24178 ? _T_27040 : 8'h0; // @[Mux.scala 19:72:@10015.4]
  assign _T_27049 = {_T_26818,_T_26817,_T_26816,_T_26815,_T_26814,_T_26821,_T_26820,_T_26819}; // @[Mux.scala 19:72:@10022.4]
  assign _T_27051 = _T_24179 ? _T_27049 : 8'h0; // @[Mux.scala 19:72:@10023.4]
  assign _T_27058 = {_T_26857,_T_26856,_T_26855,_T_26854,_T_26861,_T_26860,_T_26859,_T_26858}; // @[Mux.scala 19:72:@10030.4]
  assign _T_27060 = _T_24180 ? _T_27058 : 8'h0; // @[Mux.scala 19:72:@10031.4]
  assign _T_27067 = {_T_26896,_T_26895,_T_26894,_T_26901,_T_26900,_T_26899,_T_26898,_T_26897}; // @[Mux.scala 19:72:@10038.4]
  assign _T_27069 = _T_24181 ? _T_27067 : 8'h0; // @[Mux.scala 19:72:@10039.4]
  assign _T_27076 = {_T_26935,_T_26934,_T_26941,_T_26940,_T_26939,_T_26938,_T_26937,_T_26936}; // @[Mux.scala 19:72:@10046.4]
  assign _T_27078 = _T_24182 ? _T_27076 : 8'h0; // @[Mux.scala 19:72:@10047.4]
  assign _T_27085 = {_T_26974,_T_26981,_T_26980,_T_26979,_T_26978,_T_26977,_T_26976,_T_26975}; // @[Mux.scala 19:72:@10054.4]
  assign _T_27087 = _T_24183 ? _T_27085 : 8'h0; // @[Mux.scala 19:72:@10055.4]
  assign _T_27088 = _T_27024 | _T_27033; // @[Mux.scala 19:72:@10056.4]
  assign _T_27089 = _T_27088 | _T_27042; // @[Mux.scala 19:72:@10057.4]
  assign _T_27090 = _T_27089 | _T_27051; // @[Mux.scala 19:72:@10058.4]
  assign _T_27091 = _T_27090 | _T_27060; // @[Mux.scala 19:72:@10059.4]
  assign _T_27092 = _T_27091 | _T_27069; // @[Mux.scala 19:72:@10060.4]
  assign _T_27093 = _T_27092 | _T_27078; // @[Mux.scala 19:72:@10061.4]
  assign _T_27094 = _T_27093 | _T_27087; // @[Mux.scala 19:72:@10062.4]
  assign outputPriorityPorts_0_0 = _T_27094[0]; // @[Mux.scala 19:72:@10066.4]
  assign outputPriorityPorts_0_1 = _T_27094[1]; // @[Mux.scala 19:72:@10068.4]
  assign outputPriorityPorts_0_2 = _T_27094[2]; // @[Mux.scala 19:72:@10070.4]
  assign outputPriorityPorts_0_3 = _T_27094[3]; // @[Mux.scala 19:72:@10072.4]
  assign outputPriorityPorts_0_4 = _T_27094[4]; // @[Mux.scala 19:72:@10074.4]
  assign outputPriorityPorts_0_5 = _T_27094[5]; // @[Mux.scala 19:72:@10076.4]
  assign outputPriorityPorts_0_6 = _T_27094[6]; // @[Mux.scala 19:72:@10078.4]
  assign outputPriorityPorts_0_7 = _T_27094[7]; // @[Mux.scala 19:72:@10080.4]
  assign _T_27174 = entriesPorts_1_0 & _T_26091; // @[LoadQueue.scala 298:83:@10091.4]
  assign _T_27177 = entriesPorts_1_1 & _T_26094; // @[LoadQueue.scala 298:83:@10093.4]
  assign _T_27180 = entriesPorts_1_2 & _T_26097; // @[LoadQueue.scala 298:83:@10095.4]
  assign _T_27183 = entriesPorts_1_3 & _T_26100; // @[LoadQueue.scala 298:83:@10097.4]
  assign _T_27186 = entriesPorts_1_4 & _T_26103; // @[LoadQueue.scala 298:83:@10099.4]
  assign _T_27189 = entriesPorts_1_5 & _T_26106; // @[LoadQueue.scala 298:83:@10101.4]
  assign _T_27192 = entriesPorts_1_6 & _T_26109; // @[LoadQueue.scala 298:83:@10103.4]
  assign _T_27195 = entriesPorts_1_7 & _T_26112; // @[LoadQueue.scala 298:83:@10105.4]
  assign _T_27246 = _T_27195 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10135.4]
  assign _T_27247 = _T_27192 ? 8'h40 : _T_27246; // @[Mux.scala 31:69:@10136.4]
  assign _T_27248 = _T_27189 ? 8'h20 : _T_27247; // @[Mux.scala 31:69:@10137.4]
  assign _T_27249 = _T_27186 ? 8'h10 : _T_27248; // @[Mux.scala 31:69:@10138.4]
  assign _T_27250 = _T_27183 ? 8'h8 : _T_27249; // @[Mux.scala 31:69:@10139.4]
  assign _T_27251 = _T_27180 ? 8'h4 : _T_27250; // @[Mux.scala 31:69:@10140.4]
  assign _T_27252 = _T_27177 ? 8'h2 : _T_27251; // @[Mux.scala 31:69:@10141.4]
  assign _T_27253 = _T_27174 ? 8'h1 : _T_27252; // @[Mux.scala 31:69:@10142.4]
  assign _T_27254 = _T_27253[0]; // @[OneHot.scala 66:30:@10143.4]
  assign _T_27255 = _T_27253[1]; // @[OneHot.scala 66:30:@10144.4]
  assign _T_27256 = _T_27253[2]; // @[OneHot.scala 66:30:@10145.4]
  assign _T_27257 = _T_27253[3]; // @[OneHot.scala 66:30:@10146.4]
  assign _T_27258 = _T_27253[4]; // @[OneHot.scala 66:30:@10147.4]
  assign _T_27259 = _T_27253[5]; // @[OneHot.scala 66:30:@10148.4]
  assign _T_27260 = _T_27253[6]; // @[OneHot.scala 66:30:@10149.4]
  assign _T_27261 = _T_27253[7]; // @[OneHot.scala 66:30:@10150.4]
  assign _T_27286 = _T_27174 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10160.4]
  assign _T_27287 = _T_27195 ? 8'h40 : _T_27286; // @[Mux.scala 31:69:@10161.4]
  assign _T_27288 = _T_27192 ? 8'h20 : _T_27287; // @[Mux.scala 31:69:@10162.4]
  assign _T_27289 = _T_27189 ? 8'h10 : _T_27288; // @[Mux.scala 31:69:@10163.4]
  assign _T_27290 = _T_27186 ? 8'h8 : _T_27289; // @[Mux.scala 31:69:@10164.4]
  assign _T_27291 = _T_27183 ? 8'h4 : _T_27290; // @[Mux.scala 31:69:@10165.4]
  assign _T_27292 = _T_27180 ? 8'h2 : _T_27291; // @[Mux.scala 31:69:@10166.4]
  assign _T_27293 = _T_27177 ? 8'h1 : _T_27292; // @[Mux.scala 31:69:@10167.4]
  assign _T_27294 = _T_27293[0]; // @[OneHot.scala 66:30:@10168.4]
  assign _T_27295 = _T_27293[1]; // @[OneHot.scala 66:30:@10169.4]
  assign _T_27296 = _T_27293[2]; // @[OneHot.scala 66:30:@10170.4]
  assign _T_27297 = _T_27293[3]; // @[OneHot.scala 66:30:@10171.4]
  assign _T_27298 = _T_27293[4]; // @[OneHot.scala 66:30:@10172.4]
  assign _T_27299 = _T_27293[5]; // @[OneHot.scala 66:30:@10173.4]
  assign _T_27300 = _T_27293[6]; // @[OneHot.scala 66:30:@10174.4]
  assign _T_27301 = _T_27293[7]; // @[OneHot.scala 66:30:@10175.4]
  assign _T_27326 = _T_27177 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10185.4]
  assign _T_27327 = _T_27174 ? 8'h40 : _T_27326; // @[Mux.scala 31:69:@10186.4]
  assign _T_27328 = _T_27195 ? 8'h20 : _T_27327; // @[Mux.scala 31:69:@10187.4]
  assign _T_27329 = _T_27192 ? 8'h10 : _T_27328; // @[Mux.scala 31:69:@10188.4]
  assign _T_27330 = _T_27189 ? 8'h8 : _T_27329; // @[Mux.scala 31:69:@10189.4]
  assign _T_27331 = _T_27186 ? 8'h4 : _T_27330; // @[Mux.scala 31:69:@10190.4]
  assign _T_27332 = _T_27183 ? 8'h2 : _T_27331; // @[Mux.scala 31:69:@10191.4]
  assign _T_27333 = _T_27180 ? 8'h1 : _T_27332; // @[Mux.scala 31:69:@10192.4]
  assign _T_27334 = _T_27333[0]; // @[OneHot.scala 66:30:@10193.4]
  assign _T_27335 = _T_27333[1]; // @[OneHot.scala 66:30:@10194.4]
  assign _T_27336 = _T_27333[2]; // @[OneHot.scala 66:30:@10195.4]
  assign _T_27337 = _T_27333[3]; // @[OneHot.scala 66:30:@10196.4]
  assign _T_27338 = _T_27333[4]; // @[OneHot.scala 66:30:@10197.4]
  assign _T_27339 = _T_27333[5]; // @[OneHot.scala 66:30:@10198.4]
  assign _T_27340 = _T_27333[6]; // @[OneHot.scala 66:30:@10199.4]
  assign _T_27341 = _T_27333[7]; // @[OneHot.scala 66:30:@10200.4]
  assign _T_27366 = _T_27180 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10210.4]
  assign _T_27367 = _T_27177 ? 8'h40 : _T_27366; // @[Mux.scala 31:69:@10211.4]
  assign _T_27368 = _T_27174 ? 8'h20 : _T_27367; // @[Mux.scala 31:69:@10212.4]
  assign _T_27369 = _T_27195 ? 8'h10 : _T_27368; // @[Mux.scala 31:69:@10213.4]
  assign _T_27370 = _T_27192 ? 8'h8 : _T_27369; // @[Mux.scala 31:69:@10214.4]
  assign _T_27371 = _T_27189 ? 8'h4 : _T_27370; // @[Mux.scala 31:69:@10215.4]
  assign _T_27372 = _T_27186 ? 8'h2 : _T_27371; // @[Mux.scala 31:69:@10216.4]
  assign _T_27373 = _T_27183 ? 8'h1 : _T_27372; // @[Mux.scala 31:69:@10217.4]
  assign _T_27374 = _T_27373[0]; // @[OneHot.scala 66:30:@10218.4]
  assign _T_27375 = _T_27373[1]; // @[OneHot.scala 66:30:@10219.4]
  assign _T_27376 = _T_27373[2]; // @[OneHot.scala 66:30:@10220.4]
  assign _T_27377 = _T_27373[3]; // @[OneHot.scala 66:30:@10221.4]
  assign _T_27378 = _T_27373[4]; // @[OneHot.scala 66:30:@10222.4]
  assign _T_27379 = _T_27373[5]; // @[OneHot.scala 66:30:@10223.4]
  assign _T_27380 = _T_27373[6]; // @[OneHot.scala 66:30:@10224.4]
  assign _T_27381 = _T_27373[7]; // @[OneHot.scala 66:30:@10225.4]
  assign _T_27406 = _T_27183 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10235.4]
  assign _T_27407 = _T_27180 ? 8'h40 : _T_27406; // @[Mux.scala 31:69:@10236.4]
  assign _T_27408 = _T_27177 ? 8'h20 : _T_27407; // @[Mux.scala 31:69:@10237.4]
  assign _T_27409 = _T_27174 ? 8'h10 : _T_27408; // @[Mux.scala 31:69:@10238.4]
  assign _T_27410 = _T_27195 ? 8'h8 : _T_27409; // @[Mux.scala 31:69:@10239.4]
  assign _T_27411 = _T_27192 ? 8'h4 : _T_27410; // @[Mux.scala 31:69:@10240.4]
  assign _T_27412 = _T_27189 ? 8'h2 : _T_27411; // @[Mux.scala 31:69:@10241.4]
  assign _T_27413 = _T_27186 ? 8'h1 : _T_27412; // @[Mux.scala 31:69:@10242.4]
  assign _T_27414 = _T_27413[0]; // @[OneHot.scala 66:30:@10243.4]
  assign _T_27415 = _T_27413[1]; // @[OneHot.scala 66:30:@10244.4]
  assign _T_27416 = _T_27413[2]; // @[OneHot.scala 66:30:@10245.4]
  assign _T_27417 = _T_27413[3]; // @[OneHot.scala 66:30:@10246.4]
  assign _T_27418 = _T_27413[4]; // @[OneHot.scala 66:30:@10247.4]
  assign _T_27419 = _T_27413[5]; // @[OneHot.scala 66:30:@10248.4]
  assign _T_27420 = _T_27413[6]; // @[OneHot.scala 66:30:@10249.4]
  assign _T_27421 = _T_27413[7]; // @[OneHot.scala 66:30:@10250.4]
  assign _T_27446 = _T_27186 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10260.4]
  assign _T_27447 = _T_27183 ? 8'h40 : _T_27446; // @[Mux.scala 31:69:@10261.4]
  assign _T_27448 = _T_27180 ? 8'h20 : _T_27447; // @[Mux.scala 31:69:@10262.4]
  assign _T_27449 = _T_27177 ? 8'h10 : _T_27448; // @[Mux.scala 31:69:@10263.4]
  assign _T_27450 = _T_27174 ? 8'h8 : _T_27449; // @[Mux.scala 31:69:@10264.4]
  assign _T_27451 = _T_27195 ? 8'h4 : _T_27450; // @[Mux.scala 31:69:@10265.4]
  assign _T_27452 = _T_27192 ? 8'h2 : _T_27451; // @[Mux.scala 31:69:@10266.4]
  assign _T_27453 = _T_27189 ? 8'h1 : _T_27452; // @[Mux.scala 31:69:@10267.4]
  assign _T_27454 = _T_27453[0]; // @[OneHot.scala 66:30:@10268.4]
  assign _T_27455 = _T_27453[1]; // @[OneHot.scala 66:30:@10269.4]
  assign _T_27456 = _T_27453[2]; // @[OneHot.scala 66:30:@10270.4]
  assign _T_27457 = _T_27453[3]; // @[OneHot.scala 66:30:@10271.4]
  assign _T_27458 = _T_27453[4]; // @[OneHot.scala 66:30:@10272.4]
  assign _T_27459 = _T_27453[5]; // @[OneHot.scala 66:30:@10273.4]
  assign _T_27460 = _T_27453[6]; // @[OneHot.scala 66:30:@10274.4]
  assign _T_27461 = _T_27453[7]; // @[OneHot.scala 66:30:@10275.4]
  assign _T_27486 = _T_27189 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10285.4]
  assign _T_27487 = _T_27186 ? 8'h40 : _T_27486; // @[Mux.scala 31:69:@10286.4]
  assign _T_27488 = _T_27183 ? 8'h20 : _T_27487; // @[Mux.scala 31:69:@10287.4]
  assign _T_27489 = _T_27180 ? 8'h10 : _T_27488; // @[Mux.scala 31:69:@10288.4]
  assign _T_27490 = _T_27177 ? 8'h8 : _T_27489; // @[Mux.scala 31:69:@10289.4]
  assign _T_27491 = _T_27174 ? 8'h4 : _T_27490; // @[Mux.scala 31:69:@10290.4]
  assign _T_27492 = _T_27195 ? 8'h2 : _T_27491; // @[Mux.scala 31:69:@10291.4]
  assign _T_27493 = _T_27192 ? 8'h1 : _T_27492; // @[Mux.scala 31:69:@10292.4]
  assign _T_27494 = _T_27493[0]; // @[OneHot.scala 66:30:@10293.4]
  assign _T_27495 = _T_27493[1]; // @[OneHot.scala 66:30:@10294.4]
  assign _T_27496 = _T_27493[2]; // @[OneHot.scala 66:30:@10295.4]
  assign _T_27497 = _T_27493[3]; // @[OneHot.scala 66:30:@10296.4]
  assign _T_27498 = _T_27493[4]; // @[OneHot.scala 66:30:@10297.4]
  assign _T_27499 = _T_27493[5]; // @[OneHot.scala 66:30:@10298.4]
  assign _T_27500 = _T_27493[6]; // @[OneHot.scala 66:30:@10299.4]
  assign _T_27501 = _T_27493[7]; // @[OneHot.scala 66:30:@10300.4]
  assign _T_27526 = _T_27192 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10310.4]
  assign _T_27527 = _T_27189 ? 8'h40 : _T_27526; // @[Mux.scala 31:69:@10311.4]
  assign _T_27528 = _T_27186 ? 8'h20 : _T_27527; // @[Mux.scala 31:69:@10312.4]
  assign _T_27529 = _T_27183 ? 8'h10 : _T_27528; // @[Mux.scala 31:69:@10313.4]
  assign _T_27530 = _T_27180 ? 8'h8 : _T_27529; // @[Mux.scala 31:69:@10314.4]
  assign _T_27531 = _T_27177 ? 8'h4 : _T_27530; // @[Mux.scala 31:69:@10315.4]
  assign _T_27532 = _T_27174 ? 8'h2 : _T_27531; // @[Mux.scala 31:69:@10316.4]
  assign _T_27533 = _T_27195 ? 8'h1 : _T_27532; // @[Mux.scala 31:69:@10317.4]
  assign _T_27534 = _T_27533[0]; // @[OneHot.scala 66:30:@10318.4]
  assign _T_27535 = _T_27533[1]; // @[OneHot.scala 66:30:@10319.4]
  assign _T_27536 = _T_27533[2]; // @[OneHot.scala 66:30:@10320.4]
  assign _T_27537 = _T_27533[3]; // @[OneHot.scala 66:30:@10321.4]
  assign _T_27538 = _T_27533[4]; // @[OneHot.scala 66:30:@10322.4]
  assign _T_27539 = _T_27533[5]; // @[OneHot.scala 66:30:@10323.4]
  assign _T_27540 = _T_27533[6]; // @[OneHot.scala 66:30:@10324.4]
  assign _T_27541 = _T_27533[7]; // @[OneHot.scala 66:30:@10325.4]
  assign _T_27582 = {_T_27261,_T_27260,_T_27259,_T_27258,_T_27257,_T_27256,_T_27255,_T_27254}; // @[Mux.scala 19:72:@10341.4]
  assign _T_27584 = _T_24176 ? _T_27582 : 8'h0; // @[Mux.scala 19:72:@10342.4]
  assign _T_27591 = {_T_27300,_T_27299,_T_27298,_T_27297,_T_27296,_T_27295,_T_27294,_T_27301}; // @[Mux.scala 19:72:@10349.4]
  assign _T_27593 = _T_24177 ? _T_27591 : 8'h0; // @[Mux.scala 19:72:@10350.4]
  assign _T_27600 = {_T_27339,_T_27338,_T_27337,_T_27336,_T_27335,_T_27334,_T_27341,_T_27340}; // @[Mux.scala 19:72:@10357.4]
  assign _T_27602 = _T_24178 ? _T_27600 : 8'h0; // @[Mux.scala 19:72:@10358.4]
  assign _T_27609 = {_T_27378,_T_27377,_T_27376,_T_27375,_T_27374,_T_27381,_T_27380,_T_27379}; // @[Mux.scala 19:72:@10365.4]
  assign _T_27611 = _T_24179 ? _T_27609 : 8'h0; // @[Mux.scala 19:72:@10366.4]
  assign _T_27618 = {_T_27417,_T_27416,_T_27415,_T_27414,_T_27421,_T_27420,_T_27419,_T_27418}; // @[Mux.scala 19:72:@10373.4]
  assign _T_27620 = _T_24180 ? _T_27618 : 8'h0; // @[Mux.scala 19:72:@10374.4]
  assign _T_27627 = {_T_27456,_T_27455,_T_27454,_T_27461,_T_27460,_T_27459,_T_27458,_T_27457}; // @[Mux.scala 19:72:@10381.4]
  assign _T_27629 = _T_24181 ? _T_27627 : 8'h0; // @[Mux.scala 19:72:@10382.4]
  assign _T_27636 = {_T_27495,_T_27494,_T_27501,_T_27500,_T_27499,_T_27498,_T_27497,_T_27496}; // @[Mux.scala 19:72:@10389.4]
  assign _T_27638 = _T_24182 ? _T_27636 : 8'h0; // @[Mux.scala 19:72:@10390.4]
  assign _T_27645 = {_T_27534,_T_27541,_T_27540,_T_27539,_T_27538,_T_27537,_T_27536,_T_27535}; // @[Mux.scala 19:72:@10397.4]
  assign _T_27647 = _T_24183 ? _T_27645 : 8'h0; // @[Mux.scala 19:72:@10398.4]
  assign _T_27648 = _T_27584 | _T_27593; // @[Mux.scala 19:72:@10399.4]
  assign _T_27649 = _T_27648 | _T_27602; // @[Mux.scala 19:72:@10400.4]
  assign _T_27650 = _T_27649 | _T_27611; // @[Mux.scala 19:72:@10401.4]
  assign _T_27651 = _T_27650 | _T_27620; // @[Mux.scala 19:72:@10402.4]
  assign _T_27652 = _T_27651 | _T_27629; // @[Mux.scala 19:72:@10403.4]
  assign _T_27653 = _T_27652 | _T_27638; // @[Mux.scala 19:72:@10404.4]
  assign _T_27654 = _T_27653 | _T_27647; // @[Mux.scala 19:72:@10405.4]
  assign inputPriorityPorts_1_0 = _T_27654[0]; // @[Mux.scala 19:72:@10409.4]
  assign inputPriorityPorts_1_1 = _T_27654[1]; // @[Mux.scala 19:72:@10411.4]
  assign inputPriorityPorts_1_2 = _T_27654[2]; // @[Mux.scala 19:72:@10413.4]
  assign inputPriorityPorts_1_3 = _T_27654[3]; // @[Mux.scala 19:72:@10415.4]
  assign inputPriorityPorts_1_4 = _T_27654[4]; // @[Mux.scala 19:72:@10417.4]
  assign inputPriorityPorts_1_5 = _T_27654[5]; // @[Mux.scala 19:72:@10419.4]
  assign inputPriorityPorts_1_6 = _T_27654[6]; // @[Mux.scala 19:72:@10421.4]
  assign inputPriorityPorts_1_7 = _T_27654[7]; // @[Mux.scala 19:72:@10423.4]
  assign _T_27768 = entriesPorts_1_7 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10453.4]
  assign _T_27769 = entriesPorts_1_6 ? 8'h40 : _T_27768; // @[Mux.scala 31:69:@10454.4]
  assign _T_27770 = entriesPorts_1_5 ? 8'h20 : _T_27769; // @[Mux.scala 31:69:@10455.4]
  assign _T_27771 = entriesPorts_1_4 ? 8'h10 : _T_27770; // @[Mux.scala 31:69:@10456.4]
  assign _T_27772 = entriesPorts_1_3 ? 8'h8 : _T_27771; // @[Mux.scala 31:69:@10457.4]
  assign _T_27773 = entriesPorts_1_2 ? 8'h4 : _T_27772; // @[Mux.scala 31:69:@10458.4]
  assign _T_27774 = entriesPorts_1_1 ? 8'h2 : _T_27773; // @[Mux.scala 31:69:@10459.4]
  assign _T_27775 = entriesPorts_1_0 ? 8'h1 : _T_27774; // @[Mux.scala 31:69:@10460.4]
  assign _T_27776 = _T_27775[0]; // @[OneHot.scala 66:30:@10461.4]
  assign _T_27777 = _T_27775[1]; // @[OneHot.scala 66:30:@10462.4]
  assign _T_27778 = _T_27775[2]; // @[OneHot.scala 66:30:@10463.4]
  assign _T_27779 = _T_27775[3]; // @[OneHot.scala 66:30:@10464.4]
  assign _T_27780 = _T_27775[4]; // @[OneHot.scala 66:30:@10465.4]
  assign _T_27781 = _T_27775[5]; // @[OneHot.scala 66:30:@10466.4]
  assign _T_27782 = _T_27775[6]; // @[OneHot.scala 66:30:@10467.4]
  assign _T_27783 = _T_27775[7]; // @[OneHot.scala 66:30:@10468.4]
  assign _T_27808 = entriesPorts_1_0 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10478.4]
  assign _T_27809 = entriesPorts_1_7 ? 8'h40 : _T_27808; // @[Mux.scala 31:69:@10479.4]
  assign _T_27810 = entriesPorts_1_6 ? 8'h20 : _T_27809; // @[Mux.scala 31:69:@10480.4]
  assign _T_27811 = entriesPorts_1_5 ? 8'h10 : _T_27810; // @[Mux.scala 31:69:@10481.4]
  assign _T_27812 = entriesPorts_1_4 ? 8'h8 : _T_27811; // @[Mux.scala 31:69:@10482.4]
  assign _T_27813 = entriesPorts_1_3 ? 8'h4 : _T_27812; // @[Mux.scala 31:69:@10483.4]
  assign _T_27814 = entriesPorts_1_2 ? 8'h2 : _T_27813; // @[Mux.scala 31:69:@10484.4]
  assign _T_27815 = entriesPorts_1_1 ? 8'h1 : _T_27814; // @[Mux.scala 31:69:@10485.4]
  assign _T_27816 = _T_27815[0]; // @[OneHot.scala 66:30:@10486.4]
  assign _T_27817 = _T_27815[1]; // @[OneHot.scala 66:30:@10487.4]
  assign _T_27818 = _T_27815[2]; // @[OneHot.scala 66:30:@10488.4]
  assign _T_27819 = _T_27815[3]; // @[OneHot.scala 66:30:@10489.4]
  assign _T_27820 = _T_27815[4]; // @[OneHot.scala 66:30:@10490.4]
  assign _T_27821 = _T_27815[5]; // @[OneHot.scala 66:30:@10491.4]
  assign _T_27822 = _T_27815[6]; // @[OneHot.scala 66:30:@10492.4]
  assign _T_27823 = _T_27815[7]; // @[OneHot.scala 66:30:@10493.4]
  assign _T_27848 = entriesPorts_1_1 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10503.4]
  assign _T_27849 = entriesPorts_1_0 ? 8'h40 : _T_27848; // @[Mux.scala 31:69:@10504.4]
  assign _T_27850 = entriesPorts_1_7 ? 8'h20 : _T_27849; // @[Mux.scala 31:69:@10505.4]
  assign _T_27851 = entriesPorts_1_6 ? 8'h10 : _T_27850; // @[Mux.scala 31:69:@10506.4]
  assign _T_27852 = entriesPorts_1_5 ? 8'h8 : _T_27851; // @[Mux.scala 31:69:@10507.4]
  assign _T_27853 = entriesPorts_1_4 ? 8'h4 : _T_27852; // @[Mux.scala 31:69:@10508.4]
  assign _T_27854 = entriesPorts_1_3 ? 8'h2 : _T_27853; // @[Mux.scala 31:69:@10509.4]
  assign _T_27855 = entriesPorts_1_2 ? 8'h1 : _T_27854; // @[Mux.scala 31:69:@10510.4]
  assign _T_27856 = _T_27855[0]; // @[OneHot.scala 66:30:@10511.4]
  assign _T_27857 = _T_27855[1]; // @[OneHot.scala 66:30:@10512.4]
  assign _T_27858 = _T_27855[2]; // @[OneHot.scala 66:30:@10513.4]
  assign _T_27859 = _T_27855[3]; // @[OneHot.scala 66:30:@10514.4]
  assign _T_27860 = _T_27855[4]; // @[OneHot.scala 66:30:@10515.4]
  assign _T_27861 = _T_27855[5]; // @[OneHot.scala 66:30:@10516.4]
  assign _T_27862 = _T_27855[6]; // @[OneHot.scala 66:30:@10517.4]
  assign _T_27863 = _T_27855[7]; // @[OneHot.scala 66:30:@10518.4]
  assign _T_27888 = entriesPorts_1_2 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10528.4]
  assign _T_27889 = entriesPorts_1_1 ? 8'h40 : _T_27888; // @[Mux.scala 31:69:@10529.4]
  assign _T_27890 = entriesPorts_1_0 ? 8'h20 : _T_27889; // @[Mux.scala 31:69:@10530.4]
  assign _T_27891 = entriesPorts_1_7 ? 8'h10 : _T_27890; // @[Mux.scala 31:69:@10531.4]
  assign _T_27892 = entriesPorts_1_6 ? 8'h8 : _T_27891; // @[Mux.scala 31:69:@10532.4]
  assign _T_27893 = entriesPorts_1_5 ? 8'h4 : _T_27892; // @[Mux.scala 31:69:@10533.4]
  assign _T_27894 = entriesPorts_1_4 ? 8'h2 : _T_27893; // @[Mux.scala 31:69:@10534.4]
  assign _T_27895 = entriesPorts_1_3 ? 8'h1 : _T_27894; // @[Mux.scala 31:69:@10535.4]
  assign _T_27896 = _T_27895[0]; // @[OneHot.scala 66:30:@10536.4]
  assign _T_27897 = _T_27895[1]; // @[OneHot.scala 66:30:@10537.4]
  assign _T_27898 = _T_27895[2]; // @[OneHot.scala 66:30:@10538.4]
  assign _T_27899 = _T_27895[3]; // @[OneHot.scala 66:30:@10539.4]
  assign _T_27900 = _T_27895[4]; // @[OneHot.scala 66:30:@10540.4]
  assign _T_27901 = _T_27895[5]; // @[OneHot.scala 66:30:@10541.4]
  assign _T_27902 = _T_27895[6]; // @[OneHot.scala 66:30:@10542.4]
  assign _T_27903 = _T_27895[7]; // @[OneHot.scala 66:30:@10543.4]
  assign _T_27928 = entriesPorts_1_3 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10553.4]
  assign _T_27929 = entriesPorts_1_2 ? 8'h40 : _T_27928; // @[Mux.scala 31:69:@10554.4]
  assign _T_27930 = entriesPorts_1_1 ? 8'h20 : _T_27929; // @[Mux.scala 31:69:@10555.4]
  assign _T_27931 = entriesPorts_1_0 ? 8'h10 : _T_27930; // @[Mux.scala 31:69:@10556.4]
  assign _T_27932 = entriesPorts_1_7 ? 8'h8 : _T_27931; // @[Mux.scala 31:69:@10557.4]
  assign _T_27933 = entriesPorts_1_6 ? 8'h4 : _T_27932; // @[Mux.scala 31:69:@10558.4]
  assign _T_27934 = entriesPorts_1_5 ? 8'h2 : _T_27933; // @[Mux.scala 31:69:@10559.4]
  assign _T_27935 = entriesPorts_1_4 ? 8'h1 : _T_27934; // @[Mux.scala 31:69:@10560.4]
  assign _T_27936 = _T_27935[0]; // @[OneHot.scala 66:30:@10561.4]
  assign _T_27937 = _T_27935[1]; // @[OneHot.scala 66:30:@10562.4]
  assign _T_27938 = _T_27935[2]; // @[OneHot.scala 66:30:@10563.4]
  assign _T_27939 = _T_27935[3]; // @[OneHot.scala 66:30:@10564.4]
  assign _T_27940 = _T_27935[4]; // @[OneHot.scala 66:30:@10565.4]
  assign _T_27941 = _T_27935[5]; // @[OneHot.scala 66:30:@10566.4]
  assign _T_27942 = _T_27935[6]; // @[OneHot.scala 66:30:@10567.4]
  assign _T_27943 = _T_27935[7]; // @[OneHot.scala 66:30:@10568.4]
  assign _T_27968 = entriesPorts_1_4 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10578.4]
  assign _T_27969 = entriesPorts_1_3 ? 8'h40 : _T_27968; // @[Mux.scala 31:69:@10579.4]
  assign _T_27970 = entriesPorts_1_2 ? 8'h20 : _T_27969; // @[Mux.scala 31:69:@10580.4]
  assign _T_27971 = entriesPorts_1_1 ? 8'h10 : _T_27970; // @[Mux.scala 31:69:@10581.4]
  assign _T_27972 = entriesPorts_1_0 ? 8'h8 : _T_27971; // @[Mux.scala 31:69:@10582.4]
  assign _T_27973 = entriesPorts_1_7 ? 8'h4 : _T_27972; // @[Mux.scala 31:69:@10583.4]
  assign _T_27974 = entriesPorts_1_6 ? 8'h2 : _T_27973; // @[Mux.scala 31:69:@10584.4]
  assign _T_27975 = entriesPorts_1_5 ? 8'h1 : _T_27974; // @[Mux.scala 31:69:@10585.4]
  assign _T_27976 = _T_27975[0]; // @[OneHot.scala 66:30:@10586.4]
  assign _T_27977 = _T_27975[1]; // @[OneHot.scala 66:30:@10587.4]
  assign _T_27978 = _T_27975[2]; // @[OneHot.scala 66:30:@10588.4]
  assign _T_27979 = _T_27975[3]; // @[OneHot.scala 66:30:@10589.4]
  assign _T_27980 = _T_27975[4]; // @[OneHot.scala 66:30:@10590.4]
  assign _T_27981 = _T_27975[5]; // @[OneHot.scala 66:30:@10591.4]
  assign _T_27982 = _T_27975[6]; // @[OneHot.scala 66:30:@10592.4]
  assign _T_27983 = _T_27975[7]; // @[OneHot.scala 66:30:@10593.4]
  assign _T_28008 = entriesPorts_1_5 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10603.4]
  assign _T_28009 = entriesPorts_1_4 ? 8'h40 : _T_28008; // @[Mux.scala 31:69:@10604.4]
  assign _T_28010 = entriesPorts_1_3 ? 8'h20 : _T_28009; // @[Mux.scala 31:69:@10605.4]
  assign _T_28011 = entriesPorts_1_2 ? 8'h10 : _T_28010; // @[Mux.scala 31:69:@10606.4]
  assign _T_28012 = entriesPorts_1_1 ? 8'h8 : _T_28011; // @[Mux.scala 31:69:@10607.4]
  assign _T_28013 = entriesPorts_1_0 ? 8'h4 : _T_28012; // @[Mux.scala 31:69:@10608.4]
  assign _T_28014 = entriesPorts_1_7 ? 8'h2 : _T_28013; // @[Mux.scala 31:69:@10609.4]
  assign _T_28015 = entriesPorts_1_6 ? 8'h1 : _T_28014; // @[Mux.scala 31:69:@10610.4]
  assign _T_28016 = _T_28015[0]; // @[OneHot.scala 66:30:@10611.4]
  assign _T_28017 = _T_28015[1]; // @[OneHot.scala 66:30:@10612.4]
  assign _T_28018 = _T_28015[2]; // @[OneHot.scala 66:30:@10613.4]
  assign _T_28019 = _T_28015[3]; // @[OneHot.scala 66:30:@10614.4]
  assign _T_28020 = _T_28015[4]; // @[OneHot.scala 66:30:@10615.4]
  assign _T_28021 = _T_28015[5]; // @[OneHot.scala 66:30:@10616.4]
  assign _T_28022 = _T_28015[6]; // @[OneHot.scala 66:30:@10617.4]
  assign _T_28023 = _T_28015[7]; // @[OneHot.scala 66:30:@10618.4]
  assign _T_28048 = entriesPorts_1_6 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10628.4]
  assign _T_28049 = entriesPorts_1_5 ? 8'h40 : _T_28048; // @[Mux.scala 31:69:@10629.4]
  assign _T_28050 = entriesPorts_1_4 ? 8'h20 : _T_28049; // @[Mux.scala 31:69:@10630.4]
  assign _T_28051 = entriesPorts_1_3 ? 8'h10 : _T_28050; // @[Mux.scala 31:69:@10631.4]
  assign _T_28052 = entriesPorts_1_2 ? 8'h8 : _T_28051; // @[Mux.scala 31:69:@10632.4]
  assign _T_28053 = entriesPorts_1_1 ? 8'h4 : _T_28052; // @[Mux.scala 31:69:@10633.4]
  assign _T_28054 = entriesPorts_1_0 ? 8'h2 : _T_28053; // @[Mux.scala 31:69:@10634.4]
  assign _T_28055 = entriesPorts_1_7 ? 8'h1 : _T_28054; // @[Mux.scala 31:69:@10635.4]
  assign _T_28056 = _T_28055[0]; // @[OneHot.scala 66:30:@10636.4]
  assign _T_28057 = _T_28055[1]; // @[OneHot.scala 66:30:@10637.4]
  assign _T_28058 = _T_28055[2]; // @[OneHot.scala 66:30:@10638.4]
  assign _T_28059 = _T_28055[3]; // @[OneHot.scala 66:30:@10639.4]
  assign _T_28060 = _T_28055[4]; // @[OneHot.scala 66:30:@10640.4]
  assign _T_28061 = _T_28055[5]; // @[OneHot.scala 66:30:@10641.4]
  assign _T_28062 = _T_28055[6]; // @[OneHot.scala 66:30:@10642.4]
  assign _T_28063 = _T_28055[7]; // @[OneHot.scala 66:30:@10643.4]
  assign _T_28104 = {_T_27783,_T_27782,_T_27781,_T_27780,_T_27779,_T_27778,_T_27777,_T_27776}; // @[Mux.scala 19:72:@10659.4]
  assign _T_28106 = _T_24176 ? _T_28104 : 8'h0; // @[Mux.scala 19:72:@10660.4]
  assign _T_28113 = {_T_27822,_T_27821,_T_27820,_T_27819,_T_27818,_T_27817,_T_27816,_T_27823}; // @[Mux.scala 19:72:@10667.4]
  assign _T_28115 = _T_24177 ? _T_28113 : 8'h0; // @[Mux.scala 19:72:@10668.4]
  assign _T_28122 = {_T_27861,_T_27860,_T_27859,_T_27858,_T_27857,_T_27856,_T_27863,_T_27862}; // @[Mux.scala 19:72:@10675.4]
  assign _T_28124 = _T_24178 ? _T_28122 : 8'h0; // @[Mux.scala 19:72:@10676.4]
  assign _T_28131 = {_T_27900,_T_27899,_T_27898,_T_27897,_T_27896,_T_27903,_T_27902,_T_27901}; // @[Mux.scala 19:72:@10683.4]
  assign _T_28133 = _T_24179 ? _T_28131 : 8'h0; // @[Mux.scala 19:72:@10684.4]
  assign _T_28140 = {_T_27939,_T_27938,_T_27937,_T_27936,_T_27943,_T_27942,_T_27941,_T_27940}; // @[Mux.scala 19:72:@10691.4]
  assign _T_28142 = _T_24180 ? _T_28140 : 8'h0; // @[Mux.scala 19:72:@10692.4]
  assign _T_28149 = {_T_27978,_T_27977,_T_27976,_T_27983,_T_27982,_T_27981,_T_27980,_T_27979}; // @[Mux.scala 19:72:@10699.4]
  assign _T_28151 = _T_24181 ? _T_28149 : 8'h0; // @[Mux.scala 19:72:@10700.4]
  assign _T_28158 = {_T_28017,_T_28016,_T_28023,_T_28022,_T_28021,_T_28020,_T_28019,_T_28018}; // @[Mux.scala 19:72:@10707.4]
  assign _T_28160 = _T_24182 ? _T_28158 : 8'h0; // @[Mux.scala 19:72:@10708.4]
  assign _T_28167 = {_T_28056,_T_28063,_T_28062,_T_28061,_T_28060,_T_28059,_T_28058,_T_28057}; // @[Mux.scala 19:72:@10715.4]
  assign _T_28169 = _T_24183 ? _T_28167 : 8'h0; // @[Mux.scala 19:72:@10716.4]
  assign _T_28170 = _T_28106 | _T_28115; // @[Mux.scala 19:72:@10717.4]
  assign _T_28171 = _T_28170 | _T_28124; // @[Mux.scala 19:72:@10718.4]
  assign _T_28172 = _T_28171 | _T_28133; // @[Mux.scala 19:72:@10719.4]
  assign _T_28173 = _T_28172 | _T_28142; // @[Mux.scala 19:72:@10720.4]
  assign _T_28174 = _T_28173 | _T_28151; // @[Mux.scala 19:72:@10721.4]
  assign _T_28175 = _T_28174 | _T_28160; // @[Mux.scala 19:72:@10722.4]
  assign _T_28176 = _T_28175 | _T_28169; // @[Mux.scala 19:72:@10723.4]
  assign outputPriorityPorts_1_0 = _T_28176[0]; // @[Mux.scala 19:72:@10727.4]
  assign outputPriorityPorts_1_1 = _T_28176[1]; // @[Mux.scala 19:72:@10729.4]
  assign outputPriorityPorts_1_2 = _T_28176[2]; // @[Mux.scala 19:72:@10731.4]
  assign outputPriorityPorts_1_3 = _T_28176[3]; // @[Mux.scala 19:72:@10733.4]
  assign outputPriorityPorts_1_4 = _T_28176[4]; // @[Mux.scala 19:72:@10735.4]
  assign outputPriorityPorts_1_5 = _T_28176[5]; // @[Mux.scala 19:72:@10737.4]
  assign outputPriorityPorts_1_6 = _T_28176[6]; // @[Mux.scala 19:72:@10739.4]
  assign outputPriorityPorts_1_7 = _T_28176[7]; // @[Mux.scala 19:72:@10741.4]
  assign _T_28256 = entriesPorts_2_0 & _T_26091; // @[LoadQueue.scala 298:83:@10752.4]
  assign _T_28259 = entriesPorts_2_1 & _T_26094; // @[LoadQueue.scala 298:83:@10754.4]
  assign _T_28262 = entriesPorts_2_2 & _T_26097; // @[LoadQueue.scala 298:83:@10756.4]
  assign _T_28265 = entriesPorts_2_3 & _T_26100; // @[LoadQueue.scala 298:83:@10758.4]
  assign _T_28268 = entriesPorts_2_4 & _T_26103; // @[LoadQueue.scala 298:83:@10760.4]
  assign _T_28271 = entriesPorts_2_5 & _T_26106; // @[LoadQueue.scala 298:83:@10762.4]
  assign _T_28274 = entriesPorts_2_6 & _T_26109; // @[LoadQueue.scala 298:83:@10764.4]
  assign _T_28277 = entriesPorts_2_7 & _T_26112; // @[LoadQueue.scala 298:83:@10766.4]
  assign _T_28328 = _T_28277 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10796.4]
  assign _T_28329 = _T_28274 ? 8'h40 : _T_28328; // @[Mux.scala 31:69:@10797.4]
  assign _T_28330 = _T_28271 ? 8'h20 : _T_28329; // @[Mux.scala 31:69:@10798.4]
  assign _T_28331 = _T_28268 ? 8'h10 : _T_28330; // @[Mux.scala 31:69:@10799.4]
  assign _T_28332 = _T_28265 ? 8'h8 : _T_28331; // @[Mux.scala 31:69:@10800.4]
  assign _T_28333 = _T_28262 ? 8'h4 : _T_28332; // @[Mux.scala 31:69:@10801.4]
  assign _T_28334 = _T_28259 ? 8'h2 : _T_28333; // @[Mux.scala 31:69:@10802.4]
  assign _T_28335 = _T_28256 ? 8'h1 : _T_28334; // @[Mux.scala 31:69:@10803.4]
  assign _T_28336 = _T_28335[0]; // @[OneHot.scala 66:30:@10804.4]
  assign _T_28337 = _T_28335[1]; // @[OneHot.scala 66:30:@10805.4]
  assign _T_28338 = _T_28335[2]; // @[OneHot.scala 66:30:@10806.4]
  assign _T_28339 = _T_28335[3]; // @[OneHot.scala 66:30:@10807.4]
  assign _T_28340 = _T_28335[4]; // @[OneHot.scala 66:30:@10808.4]
  assign _T_28341 = _T_28335[5]; // @[OneHot.scala 66:30:@10809.4]
  assign _T_28342 = _T_28335[6]; // @[OneHot.scala 66:30:@10810.4]
  assign _T_28343 = _T_28335[7]; // @[OneHot.scala 66:30:@10811.4]
  assign _T_28368 = _T_28256 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10821.4]
  assign _T_28369 = _T_28277 ? 8'h40 : _T_28368; // @[Mux.scala 31:69:@10822.4]
  assign _T_28370 = _T_28274 ? 8'h20 : _T_28369; // @[Mux.scala 31:69:@10823.4]
  assign _T_28371 = _T_28271 ? 8'h10 : _T_28370; // @[Mux.scala 31:69:@10824.4]
  assign _T_28372 = _T_28268 ? 8'h8 : _T_28371; // @[Mux.scala 31:69:@10825.4]
  assign _T_28373 = _T_28265 ? 8'h4 : _T_28372; // @[Mux.scala 31:69:@10826.4]
  assign _T_28374 = _T_28262 ? 8'h2 : _T_28373; // @[Mux.scala 31:69:@10827.4]
  assign _T_28375 = _T_28259 ? 8'h1 : _T_28374; // @[Mux.scala 31:69:@10828.4]
  assign _T_28376 = _T_28375[0]; // @[OneHot.scala 66:30:@10829.4]
  assign _T_28377 = _T_28375[1]; // @[OneHot.scala 66:30:@10830.4]
  assign _T_28378 = _T_28375[2]; // @[OneHot.scala 66:30:@10831.4]
  assign _T_28379 = _T_28375[3]; // @[OneHot.scala 66:30:@10832.4]
  assign _T_28380 = _T_28375[4]; // @[OneHot.scala 66:30:@10833.4]
  assign _T_28381 = _T_28375[5]; // @[OneHot.scala 66:30:@10834.4]
  assign _T_28382 = _T_28375[6]; // @[OneHot.scala 66:30:@10835.4]
  assign _T_28383 = _T_28375[7]; // @[OneHot.scala 66:30:@10836.4]
  assign _T_28408 = _T_28259 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10846.4]
  assign _T_28409 = _T_28256 ? 8'h40 : _T_28408; // @[Mux.scala 31:69:@10847.4]
  assign _T_28410 = _T_28277 ? 8'h20 : _T_28409; // @[Mux.scala 31:69:@10848.4]
  assign _T_28411 = _T_28274 ? 8'h10 : _T_28410; // @[Mux.scala 31:69:@10849.4]
  assign _T_28412 = _T_28271 ? 8'h8 : _T_28411; // @[Mux.scala 31:69:@10850.4]
  assign _T_28413 = _T_28268 ? 8'h4 : _T_28412; // @[Mux.scala 31:69:@10851.4]
  assign _T_28414 = _T_28265 ? 8'h2 : _T_28413; // @[Mux.scala 31:69:@10852.4]
  assign _T_28415 = _T_28262 ? 8'h1 : _T_28414; // @[Mux.scala 31:69:@10853.4]
  assign _T_28416 = _T_28415[0]; // @[OneHot.scala 66:30:@10854.4]
  assign _T_28417 = _T_28415[1]; // @[OneHot.scala 66:30:@10855.4]
  assign _T_28418 = _T_28415[2]; // @[OneHot.scala 66:30:@10856.4]
  assign _T_28419 = _T_28415[3]; // @[OneHot.scala 66:30:@10857.4]
  assign _T_28420 = _T_28415[4]; // @[OneHot.scala 66:30:@10858.4]
  assign _T_28421 = _T_28415[5]; // @[OneHot.scala 66:30:@10859.4]
  assign _T_28422 = _T_28415[6]; // @[OneHot.scala 66:30:@10860.4]
  assign _T_28423 = _T_28415[7]; // @[OneHot.scala 66:30:@10861.4]
  assign _T_28448 = _T_28262 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10871.4]
  assign _T_28449 = _T_28259 ? 8'h40 : _T_28448; // @[Mux.scala 31:69:@10872.4]
  assign _T_28450 = _T_28256 ? 8'h20 : _T_28449; // @[Mux.scala 31:69:@10873.4]
  assign _T_28451 = _T_28277 ? 8'h10 : _T_28450; // @[Mux.scala 31:69:@10874.4]
  assign _T_28452 = _T_28274 ? 8'h8 : _T_28451; // @[Mux.scala 31:69:@10875.4]
  assign _T_28453 = _T_28271 ? 8'h4 : _T_28452; // @[Mux.scala 31:69:@10876.4]
  assign _T_28454 = _T_28268 ? 8'h2 : _T_28453; // @[Mux.scala 31:69:@10877.4]
  assign _T_28455 = _T_28265 ? 8'h1 : _T_28454; // @[Mux.scala 31:69:@10878.4]
  assign _T_28456 = _T_28455[0]; // @[OneHot.scala 66:30:@10879.4]
  assign _T_28457 = _T_28455[1]; // @[OneHot.scala 66:30:@10880.4]
  assign _T_28458 = _T_28455[2]; // @[OneHot.scala 66:30:@10881.4]
  assign _T_28459 = _T_28455[3]; // @[OneHot.scala 66:30:@10882.4]
  assign _T_28460 = _T_28455[4]; // @[OneHot.scala 66:30:@10883.4]
  assign _T_28461 = _T_28455[5]; // @[OneHot.scala 66:30:@10884.4]
  assign _T_28462 = _T_28455[6]; // @[OneHot.scala 66:30:@10885.4]
  assign _T_28463 = _T_28455[7]; // @[OneHot.scala 66:30:@10886.4]
  assign _T_28488 = _T_28265 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10896.4]
  assign _T_28489 = _T_28262 ? 8'h40 : _T_28488; // @[Mux.scala 31:69:@10897.4]
  assign _T_28490 = _T_28259 ? 8'h20 : _T_28489; // @[Mux.scala 31:69:@10898.4]
  assign _T_28491 = _T_28256 ? 8'h10 : _T_28490; // @[Mux.scala 31:69:@10899.4]
  assign _T_28492 = _T_28277 ? 8'h8 : _T_28491; // @[Mux.scala 31:69:@10900.4]
  assign _T_28493 = _T_28274 ? 8'h4 : _T_28492; // @[Mux.scala 31:69:@10901.4]
  assign _T_28494 = _T_28271 ? 8'h2 : _T_28493; // @[Mux.scala 31:69:@10902.4]
  assign _T_28495 = _T_28268 ? 8'h1 : _T_28494; // @[Mux.scala 31:69:@10903.4]
  assign _T_28496 = _T_28495[0]; // @[OneHot.scala 66:30:@10904.4]
  assign _T_28497 = _T_28495[1]; // @[OneHot.scala 66:30:@10905.4]
  assign _T_28498 = _T_28495[2]; // @[OneHot.scala 66:30:@10906.4]
  assign _T_28499 = _T_28495[3]; // @[OneHot.scala 66:30:@10907.4]
  assign _T_28500 = _T_28495[4]; // @[OneHot.scala 66:30:@10908.4]
  assign _T_28501 = _T_28495[5]; // @[OneHot.scala 66:30:@10909.4]
  assign _T_28502 = _T_28495[6]; // @[OneHot.scala 66:30:@10910.4]
  assign _T_28503 = _T_28495[7]; // @[OneHot.scala 66:30:@10911.4]
  assign _T_28528 = _T_28268 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10921.4]
  assign _T_28529 = _T_28265 ? 8'h40 : _T_28528; // @[Mux.scala 31:69:@10922.4]
  assign _T_28530 = _T_28262 ? 8'h20 : _T_28529; // @[Mux.scala 31:69:@10923.4]
  assign _T_28531 = _T_28259 ? 8'h10 : _T_28530; // @[Mux.scala 31:69:@10924.4]
  assign _T_28532 = _T_28256 ? 8'h8 : _T_28531; // @[Mux.scala 31:69:@10925.4]
  assign _T_28533 = _T_28277 ? 8'h4 : _T_28532; // @[Mux.scala 31:69:@10926.4]
  assign _T_28534 = _T_28274 ? 8'h2 : _T_28533; // @[Mux.scala 31:69:@10927.4]
  assign _T_28535 = _T_28271 ? 8'h1 : _T_28534; // @[Mux.scala 31:69:@10928.4]
  assign _T_28536 = _T_28535[0]; // @[OneHot.scala 66:30:@10929.4]
  assign _T_28537 = _T_28535[1]; // @[OneHot.scala 66:30:@10930.4]
  assign _T_28538 = _T_28535[2]; // @[OneHot.scala 66:30:@10931.4]
  assign _T_28539 = _T_28535[3]; // @[OneHot.scala 66:30:@10932.4]
  assign _T_28540 = _T_28535[4]; // @[OneHot.scala 66:30:@10933.4]
  assign _T_28541 = _T_28535[5]; // @[OneHot.scala 66:30:@10934.4]
  assign _T_28542 = _T_28535[6]; // @[OneHot.scala 66:30:@10935.4]
  assign _T_28543 = _T_28535[7]; // @[OneHot.scala 66:30:@10936.4]
  assign _T_28568 = _T_28271 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10946.4]
  assign _T_28569 = _T_28268 ? 8'h40 : _T_28568; // @[Mux.scala 31:69:@10947.4]
  assign _T_28570 = _T_28265 ? 8'h20 : _T_28569; // @[Mux.scala 31:69:@10948.4]
  assign _T_28571 = _T_28262 ? 8'h10 : _T_28570; // @[Mux.scala 31:69:@10949.4]
  assign _T_28572 = _T_28259 ? 8'h8 : _T_28571; // @[Mux.scala 31:69:@10950.4]
  assign _T_28573 = _T_28256 ? 8'h4 : _T_28572; // @[Mux.scala 31:69:@10951.4]
  assign _T_28574 = _T_28277 ? 8'h2 : _T_28573; // @[Mux.scala 31:69:@10952.4]
  assign _T_28575 = _T_28274 ? 8'h1 : _T_28574; // @[Mux.scala 31:69:@10953.4]
  assign _T_28576 = _T_28575[0]; // @[OneHot.scala 66:30:@10954.4]
  assign _T_28577 = _T_28575[1]; // @[OneHot.scala 66:30:@10955.4]
  assign _T_28578 = _T_28575[2]; // @[OneHot.scala 66:30:@10956.4]
  assign _T_28579 = _T_28575[3]; // @[OneHot.scala 66:30:@10957.4]
  assign _T_28580 = _T_28575[4]; // @[OneHot.scala 66:30:@10958.4]
  assign _T_28581 = _T_28575[5]; // @[OneHot.scala 66:30:@10959.4]
  assign _T_28582 = _T_28575[6]; // @[OneHot.scala 66:30:@10960.4]
  assign _T_28583 = _T_28575[7]; // @[OneHot.scala 66:30:@10961.4]
  assign _T_28608 = _T_28274 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10971.4]
  assign _T_28609 = _T_28271 ? 8'h40 : _T_28608; // @[Mux.scala 31:69:@10972.4]
  assign _T_28610 = _T_28268 ? 8'h20 : _T_28609; // @[Mux.scala 31:69:@10973.4]
  assign _T_28611 = _T_28265 ? 8'h10 : _T_28610; // @[Mux.scala 31:69:@10974.4]
  assign _T_28612 = _T_28262 ? 8'h8 : _T_28611; // @[Mux.scala 31:69:@10975.4]
  assign _T_28613 = _T_28259 ? 8'h4 : _T_28612; // @[Mux.scala 31:69:@10976.4]
  assign _T_28614 = _T_28256 ? 8'h2 : _T_28613; // @[Mux.scala 31:69:@10977.4]
  assign _T_28615 = _T_28277 ? 8'h1 : _T_28614; // @[Mux.scala 31:69:@10978.4]
  assign _T_28616 = _T_28615[0]; // @[OneHot.scala 66:30:@10979.4]
  assign _T_28617 = _T_28615[1]; // @[OneHot.scala 66:30:@10980.4]
  assign _T_28618 = _T_28615[2]; // @[OneHot.scala 66:30:@10981.4]
  assign _T_28619 = _T_28615[3]; // @[OneHot.scala 66:30:@10982.4]
  assign _T_28620 = _T_28615[4]; // @[OneHot.scala 66:30:@10983.4]
  assign _T_28621 = _T_28615[5]; // @[OneHot.scala 66:30:@10984.4]
  assign _T_28622 = _T_28615[6]; // @[OneHot.scala 66:30:@10985.4]
  assign _T_28623 = _T_28615[7]; // @[OneHot.scala 66:30:@10986.4]
  assign _T_28664 = {_T_28343,_T_28342,_T_28341,_T_28340,_T_28339,_T_28338,_T_28337,_T_28336}; // @[Mux.scala 19:72:@11002.4]
  assign _T_28666 = _T_24176 ? _T_28664 : 8'h0; // @[Mux.scala 19:72:@11003.4]
  assign _T_28673 = {_T_28382,_T_28381,_T_28380,_T_28379,_T_28378,_T_28377,_T_28376,_T_28383}; // @[Mux.scala 19:72:@11010.4]
  assign _T_28675 = _T_24177 ? _T_28673 : 8'h0; // @[Mux.scala 19:72:@11011.4]
  assign _T_28682 = {_T_28421,_T_28420,_T_28419,_T_28418,_T_28417,_T_28416,_T_28423,_T_28422}; // @[Mux.scala 19:72:@11018.4]
  assign _T_28684 = _T_24178 ? _T_28682 : 8'h0; // @[Mux.scala 19:72:@11019.4]
  assign _T_28691 = {_T_28460,_T_28459,_T_28458,_T_28457,_T_28456,_T_28463,_T_28462,_T_28461}; // @[Mux.scala 19:72:@11026.4]
  assign _T_28693 = _T_24179 ? _T_28691 : 8'h0; // @[Mux.scala 19:72:@11027.4]
  assign _T_28700 = {_T_28499,_T_28498,_T_28497,_T_28496,_T_28503,_T_28502,_T_28501,_T_28500}; // @[Mux.scala 19:72:@11034.4]
  assign _T_28702 = _T_24180 ? _T_28700 : 8'h0; // @[Mux.scala 19:72:@11035.4]
  assign _T_28709 = {_T_28538,_T_28537,_T_28536,_T_28543,_T_28542,_T_28541,_T_28540,_T_28539}; // @[Mux.scala 19:72:@11042.4]
  assign _T_28711 = _T_24181 ? _T_28709 : 8'h0; // @[Mux.scala 19:72:@11043.4]
  assign _T_28718 = {_T_28577,_T_28576,_T_28583,_T_28582,_T_28581,_T_28580,_T_28579,_T_28578}; // @[Mux.scala 19:72:@11050.4]
  assign _T_28720 = _T_24182 ? _T_28718 : 8'h0; // @[Mux.scala 19:72:@11051.4]
  assign _T_28727 = {_T_28616,_T_28623,_T_28622,_T_28621,_T_28620,_T_28619,_T_28618,_T_28617}; // @[Mux.scala 19:72:@11058.4]
  assign _T_28729 = _T_24183 ? _T_28727 : 8'h0; // @[Mux.scala 19:72:@11059.4]
  assign _T_28730 = _T_28666 | _T_28675; // @[Mux.scala 19:72:@11060.4]
  assign _T_28731 = _T_28730 | _T_28684; // @[Mux.scala 19:72:@11061.4]
  assign _T_28732 = _T_28731 | _T_28693; // @[Mux.scala 19:72:@11062.4]
  assign _T_28733 = _T_28732 | _T_28702; // @[Mux.scala 19:72:@11063.4]
  assign _T_28734 = _T_28733 | _T_28711; // @[Mux.scala 19:72:@11064.4]
  assign _T_28735 = _T_28734 | _T_28720; // @[Mux.scala 19:72:@11065.4]
  assign _T_28736 = _T_28735 | _T_28729; // @[Mux.scala 19:72:@11066.4]
  assign inputPriorityPorts_2_0 = _T_28736[0]; // @[Mux.scala 19:72:@11070.4]
  assign inputPriorityPorts_2_1 = _T_28736[1]; // @[Mux.scala 19:72:@11072.4]
  assign inputPriorityPorts_2_2 = _T_28736[2]; // @[Mux.scala 19:72:@11074.4]
  assign inputPriorityPorts_2_3 = _T_28736[3]; // @[Mux.scala 19:72:@11076.4]
  assign inputPriorityPorts_2_4 = _T_28736[4]; // @[Mux.scala 19:72:@11078.4]
  assign inputPriorityPorts_2_5 = _T_28736[5]; // @[Mux.scala 19:72:@11080.4]
  assign inputPriorityPorts_2_6 = _T_28736[6]; // @[Mux.scala 19:72:@11082.4]
  assign inputPriorityPorts_2_7 = _T_28736[7]; // @[Mux.scala 19:72:@11084.4]
  assign _T_28850 = entriesPorts_2_7 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11114.4]
  assign _T_28851 = entriesPorts_2_6 ? 8'h40 : _T_28850; // @[Mux.scala 31:69:@11115.4]
  assign _T_28852 = entriesPorts_2_5 ? 8'h20 : _T_28851; // @[Mux.scala 31:69:@11116.4]
  assign _T_28853 = entriesPorts_2_4 ? 8'h10 : _T_28852; // @[Mux.scala 31:69:@11117.4]
  assign _T_28854 = entriesPorts_2_3 ? 8'h8 : _T_28853; // @[Mux.scala 31:69:@11118.4]
  assign _T_28855 = entriesPorts_2_2 ? 8'h4 : _T_28854; // @[Mux.scala 31:69:@11119.4]
  assign _T_28856 = entriesPorts_2_1 ? 8'h2 : _T_28855; // @[Mux.scala 31:69:@11120.4]
  assign _T_28857 = entriesPorts_2_0 ? 8'h1 : _T_28856; // @[Mux.scala 31:69:@11121.4]
  assign _T_28858 = _T_28857[0]; // @[OneHot.scala 66:30:@11122.4]
  assign _T_28859 = _T_28857[1]; // @[OneHot.scala 66:30:@11123.4]
  assign _T_28860 = _T_28857[2]; // @[OneHot.scala 66:30:@11124.4]
  assign _T_28861 = _T_28857[3]; // @[OneHot.scala 66:30:@11125.4]
  assign _T_28862 = _T_28857[4]; // @[OneHot.scala 66:30:@11126.4]
  assign _T_28863 = _T_28857[5]; // @[OneHot.scala 66:30:@11127.4]
  assign _T_28864 = _T_28857[6]; // @[OneHot.scala 66:30:@11128.4]
  assign _T_28865 = _T_28857[7]; // @[OneHot.scala 66:30:@11129.4]
  assign _T_28890 = entriesPorts_2_0 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11139.4]
  assign _T_28891 = entriesPorts_2_7 ? 8'h40 : _T_28890; // @[Mux.scala 31:69:@11140.4]
  assign _T_28892 = entriesPorts_2_6 ? 8'h20 : _T_28891; // @[Mux.scala 31:69:@11141.4]
  assign _T_28893 = entriesPorts_2_5 ? 8'h10 : _T_28892; // @[Mux.scala 31:69:@11142.4]
  assign _T_28894 = entriesPorts_2_4 ? 8'h8 : _T_28893; // @[Mux.scala 31:69:@11143.4]
  assign _T_28895 = entriesPorts_2_3 ? 8'h4 : _T_28894; // @[Mux.scala 31:69:@11144.4]
  assign _T_28896 = entriesPorts_2_2 ? 8'h2 : _T_28895; // @[Mux.scala 31:69:@11145.4]
  assign _T_28897 = entriesPorts_2_1 ? 8'h1 : _T_28896; // @[Mux.scala 31:69:@11146.4]
  assign _T_28898 = _T_28897[0]; // @[OneHot.scala 66:30:@11147.4]
  assign _T_28899 = _T_28897[1]; // @[OneHot.scala 66:30:@11148.4]
  assign _T_28900 = _T_28897[2]; // @[OneHot.scala 66:30:@11149.4]
  assign _T_28901 = _T_28897[3]; // @[OneHot.scala 66:30:@11150.4]
  assign _T_28902 = _T_28897[4]; // @[OneHot.scala 66:30:@11151.4]
  assign _T_28903 = _T_28897[5]; // @[OneHot.scala 66:30:@11152.4]
  assign _T_28904 = _T_28897[6]; // @[OneHot.scala 66:30:@11153.4]
  assign _T_28905 = _T_28897[7]; // @[OneHot.scala 66:30:@11154.4]
  assign _T_28930 = entriesPorts_2_1 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11164.4]
  assign _T_28931 = entriesPorts_2_0 ? 8'h40 : _T_28930; // @[Mux.scala 31:69:@11165.4]
  assign _T_28932 = entriesPorts_2_7 ? 8'h20 : _T_28931; // @[Mux.scala 31:69:@11166.4]
  assign _T_28933 = entriesPorts_2_6 ? 8'h10 : _T_28932; // @[Mux.scala 31:69:@11167.4]
  assign _T_28934 = entriesPorts_2_5 ? 8'h8 : _T_28933; // @[Mux.scala 31:69:@11168.4]
  assign _T_28935 = entriesPorts_2_4 ? 8'h4 : _T_28934; // @[Mux.scala 31:69:@11169.4]
  assign _T_28936 = entriesPorts_2_3 ? 8'h2 : _T_28935; // @[Mux.scala 31:69:@11170.4]
  assign _T_28937 = entriesPorts_2_2 ? 8'h1 : _T_28936; // @[Mux.scala 31:69:@11171.4]
  assign _T_28938 = _T_28937[0]; // @[OneHot.scala 66:30:@11172.4]
  assign _T_28939 = _T_28937[1]; // @[OneHot.scala 66:30:@11173.4]
  assign _T_28940 = _T_28937[2]; // @[OneHot.scala 66:30:@11174.4]
  assign _T_28941 = _T_28937[3]; // @[OneHot.scala 66:30:@11175.4]
  assign _T_28942 = _T_28937[4]; // @[OneHot.scala 66:30:@11176.4]
  assign _T_28943 = _T_28937[5]; // @[OneHot.scala 66:30:@11177.4]
  assign _T_28944 = _T_28937[6]; // @[OneHot.scala 66:30:@11178.4]
  assign _T_28945 = _T_28937[7]; // @[OneHot.scala 66:30:@11179.4]
  assign _T_28970 = entriesPorts_2_2 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11189.4]
  assign _T_28971 = entriesPorts_2_1 ? 8'h40 : _T_28970; // @[Mux.scala 31:69:@11190.4]
  assign _T_28972 = entriesPorts_2_0 ? 8'h20 : _T_28971; // @[Mux.scala 31:69:@11191.4]
  assign _T_28973 = entriesPorts_2_7 ? 8'h10 : _T_28972; // @[Mux.scala 31:69:@11192.4]
  assign _T_28974 = entriesPorts_2_6 ? 8'h8 : _T_28973; // @[Mux.scala 31:69:@11193.4]
  assign _T_28975 = entriesPorts_2_5 ? 8'h4 : _T_28974; // @[Mux.scala 31:69:@11194.4]
  assign _T_28976 = entriesPorts_2_4 ? 8'h2 : _T_28975; // @[Mux.scala 31:69:@11195.4]
  assign _T_28977 = entriesPorts_2_3 ? 8'h1 : _T_28976; // @[Mux.scala 31:69:@11196.4]
  assign _T_28978 = _T_28977[0]; // @[OneHot.scala 66:30:@11197.4]
  assign _T_28979 = _T_28977[1]; // @[OneHot.scala 66:30:@11198.4]
  assign _T_28980 = _T_28977[2]; // @[OneHot.scala 66:30:@11199.4]
  assign _T_28981 = _T_28977[3]; // @[OneHot.scala 66:30:@11200.4]
  assign _T_28982 = _T_28977[4]; // @[OneHot.scala 66:30:@11201.4]
  assign _T_28983 = _T_28977[5]; // @[OneHot.scala 66:30:@11202.4]
  assign _T_28984 = _T_28977[6]; // @[OneHot.scala 66:30:@11203.4]
  assign _T_28985 = _T_28977[7]; // @[OneHot.scala 66:30:@11204.4]
  assign _T_29010 = entriesPorts_2_3 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11214.4]
  assign _T_29011 = entriesPorts_2_2 ? 8'h40 : _T_29010; // @[Mux.scala 31:69:@11215.4]
  assign _T_29012 = entriesPorts_2_1 ? 8'h20 : _T_29011; // @[Mux.scala 31:69:@11216.4]
  assign _T_29013 = entriesPorts_2_0 ? 8'h10 : _T_29012; // @[Mux.scala 31:69:@11217.4]
  assign _T_29014 = entriesPorts_2_7 ? 8'h8 : _T_29013; // @[Mux.scala 31:69:@11218.4]
  assign _T_29015 = entriesPorts_2_6 ? 8'h4 : _T_29014; // @[Mux.scala 31:69:@11219.4]
  assign _T_29016 = entriesPorts_2_5 ? 8'h2 : _T_29015; // @[Mux.scala 31:69:@11220.4]
  assign _T_29017 = entriesPorts_2_4 ? 8'h1 : _T_29016; // @[Mux.scala 31:69:@11221.4]
  assign _T_29018 = _T_29017[0]; // @[OneHot.scala 66:30:@11222.4]
  assign _T_29019 = _T_29017[1]; // @[OneHot.scala 66:30:@11223.4]
  assign _T_29020 = _T_29017[2]; // @[OneHot.scala 66:30:@11224.4]
  assign _T_29021 = _T_29017[3]; // @[OneHot.scala 66:30:@11225.4]
  assign _T_29022 = _T_29017[4]; // @[OneHot.scala 66:30:@11226.4]
  assign _T_29023 = _T_29017[5]; // @[OneHot.scala 66:30:@11227.4]
  assign _T_29024 = _T_29017[6]; // @[OneHot.scala 66:30:@11228.4]
  assign _T_29025 = _T_29017[7]; // @[OneHot.scala 66:30:@11229.4]
  assign _T_29050 = entriesPorts_2_4 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11239.4]
  assign _T_29051 = entriesPorts_2_3 ? 8'h40 : _T_29050; // @[Mux.scala 31:69:@11240.4]
  assign _T_29052 = entriesPorts_2_2 ? 8'h20 : _T_29051; // @[Mux.scala 31:69:@11241.4]
  assign _T_29053 = entriesPorts_2_1 ? 8'h10 : _T_29052; // @[Mux.scala 31:69:@11242.4]
  assign _T_29054 = entriesPorts_2_0 ? 8'h8 : _T_29053; // @[Mux.scala 31:69:@11243.4]
  assign _T_29055 = entriesPorts_2_7 ? 8'h4 : _T_29054; // @[Mux.scala 31:69:@11244.4]
  assign _T_29056 = entriesPorts_2_6 ? 8'h2 : _T_29055; // @[Mux.scala 31:69:@11245.4]
  assign _T_29057 = entriesPorts_2_5 ? 8'h1 : _T_29056; // @[Mux.scala 31:69:@11246.4]
  assign _T_29058 = _T_29057[0]; // @[OneHot.scala 66:30:@11247.4]
  assign _T_29059 = _T_29057[1]; // @[OneHot.scala 66:30:@11248.4]
  assign _T_29060 = _T_29057[2]; // @[OneHot.scala 66:30:@11249.4]
  assign _T_29061 = _T_29057[3]; // @[OneHot.scala 66:30:@11250.4]
  assign _T_29062 = _T_29057[4]; // @[OneHot.scala 66:30:@11251.4]
  assign _T_29063 = _T_29057[5]; // @[OneHot.scala 66:30:@11252.4]
  assign _T_29064 = _T_29057[6]; // @[OneHot.scala 66:30:@11253.4]
  assign _T_29065 = _T_29057[7]; // @[OneHot.scala 66:30:@11254.4]
  assign _T_29090 = entriesPorts_2_5 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11264.4]
  assign _T_29091 = entriesPorts_2_4 ? 8'h40 : _T_29090; // @[Mux.scala 31:69:@11265.4]
  assign _T_29092 = entriesPorts_2_3 ? 8'h20 : _T_29091; // @[Mux.scala 31:69:@11266.4]
  assign _T_29093 = entriesPorts_2_2 ? 8'h10 : _T_29092; // @[Mux.scala 31:69:@11267.4]
  assign _T_29094 = entriesPorts_2_1 ? 8'h8 : _T_29093; // @[Mux.scala 31:69:@11268.4]
  assign _T_29095 = entriesPorts_2_0 ? 8'h4 : _T_29094; // @[Mux.scala 31:69:@11269.4]
  assign _T_29096 = entriesPorts_2_7 ? 8'h2 : _T_29095; // @[Mux.scala 31:69:@11270.4]
  assign _T_29097 = entriesPorts_2_6 ? 8'h1 : _T_29096; // @[Mux.scala 31:69:@11271.4]
  assign _T_29098 = _T_29097[0]; // @[OneHot.scala 66:30:@11272.4]
  assign _T_29099 = _T_29097[1]; // @[OneHot.scala 66:30:@11273.4]
  assign _T_29100 = _T_29097[2]; // @[OneHot.scala 66:30:@11274.4]
  assign _T_29101 = _T_29097[3]; // @[OneHot.scala 66:30:@11275.4]
  assign _T_29102 = _T_29097[4]; // @[OneHot.scala 66:30:@11276.4]
  assign _T_29103 = _T_29097[5]; // @[OneHot.scala 66:30:@11277.4]
  assign _T_29104 = _T_29097[6]; // @[OneHot.scala 66:30:@11278.4]
  assign _T_29105 = _T_29097[7]; // @[OneHot.scala 66:30:@11279.4]
  assign _T_29130 = entriesPorts_2_6 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11289.4]
  assign _T_29131 = entriesPorts_2_5 ? 8'h40 : _T_29130; // @[Mux.scala 31:69:@11290.4]
  assign _T_29132 = entriesPorts_2_4 ? 8'h20 : _T_29131; // @[Mux.scala 31:69:@11291.4]
  assign _T_29133 = entriesPorts_2_3 ? 8'h10 : _T_29132; // @[Mux.scala 31:69:@11292.4]
  assign _T_29134 = entriesPorts_2_2 ? 8'h8 : _T_29133; // @[Mux.scala 31:69:@11293.4]
  assign _T_29135 = entriesPorts_2_1 ? 8'h4 : _T_29134; // @[Mux.scala 31:69:@11294.4]
  assign _T_29136 = entriesPorts_2_0 ? 8'h2 : _T_29135; // @[Mux.scala 31:69:@11295.4]
  assign _T_29137 = entriesPorts_2_7 ? 8'h1 : _T_29136; // @[Mux.scala 31:69:@11296.4]
  assign _T_29138 = _T_29137[0]; // @[OneHot.scala 66:30:@11297.4]
  assign _T_29139 = _T_29137[1]; // @[OneHot.scala 66:30:@11298.4]
  assign _T_29140 = _T_29137[2]; // @[OneHot.scala 66:30:@11299.4]
  assign _T_29141 = _T_29137[3]; // @[OneHot.scala 66:30:@11300.4]
  assign _T_29142 = _T_29137[4]; // @[OneHot.scala 66:30:@11301.4]
  assign _T_29143 = _T_29137[5]; // @[OneHot.scala 66:30:@11302.4]
  assign _T_29144 = _T_29137[6]; // @[OneHot.scala 66:30:@11303.4]
  assign _T_29145 = _T_29137[7]; // @[OneHot.scala 66:30:@11304.4]
  assign _T_29186 = {_T_28865,_T_28864,_T_28863,_T_28862,_T_28861,_T_28860,_T_28859,_T_28858}; // @[Mux.scala 19:72:@11320.4]
  assign _T_29188 = _T_24176 ? _T_29186 : 8'h0; // @[Mux.scala 19:72:@11321.4]
  assign _T_29195 = {_T_28904,_T_28903,_T_28902,_T_28901,_T_28900,_T_28899,_T_28898,_T_28905}; // @[Mux.scala 19:72:@11328.4]
  assign _T_29197 = _T_24177 ? _T_29195 : 8'h0; // @[Mux.scala 19:72:@11329.4]
  assign _T_29204 = {_T_28943,_T_28942,_T_28941,_T_28940,_T_28939,_T_28938,_T_28945,_T_28944}; // @[Mux.scala 19:72:@11336.4]
  assign _T_29206 = _T_24178 ? _T_29204 : 8'h0; // @[Mux.scala 19:72:@11337.4]
  assign _T_29213 = {_T_28982,_T_28981,_T_28980,_T_28979,_T_28978,_T_28985,_T_28984,_T_28983}; // @[Mux.scala 19:72:@11344.4]
  assign _T_29215 = _T_24179 ? _T_29213 : 8'h0; // @[Mux.scala 19:72:@11345.4]
  assign _T_29222 = {_T_29021,_T_29020,_T_29019,_T_29018,_T_29025,_T_29024,_T_29023,_T_29022}; // @[Mux.scala 19:72:@11352.4]
  assign _T_29224 = _T_24180 ? _T_29222 : 8'h0; // @[Mux.scala 19:72:@11353.4]
  assign _T_29231 = {_T_29060,_T_29059,_T_29058,_T_29065,_T_29064,_T_29063,_T_29062,_T_29061}; // @[Mux.scala 19:72:@11360.4]
  assign _T_29233 = _T_24181 ? _T_29231 : 8'h0; // @[Mux.scala 19:72:@11361.4]
  assign _T_29240 = {_T_29099,_T_29098,_T_29105,_T_29104,_T_29103,_T_29102,_T_29101,_T_29100}; // @[Mux.scala 19:72:@11368.4]
  assign _T_29242 = _T_24182 ? _T_29240 : 8'h0; // @[Mux.scala 19:72:@11369.4]
  assign _T_29249 = {_T_29138,_T_29145,_T_29144,_T_29143,_T_29142,_T_29141,_T_29140,_T_29139}; // @[Mux.scala 19:72:@11376.4]
  assign _T_29251 = _T_24183 ? _T_29249 : 8'h0; // @[Mux.scala 19:72:@11377.4]
  assign _T_29252 = _T_29188 | _T_29197; // @[Mux.scala 19:72:@11378.4]
  assign _T_29253 = _T_29252 | _T_29206; // @[Mux.scala 19:72:@11379.4]
  assign _T_29254 = _T_29253 | _T_29215; // @[Mux.scala 19:72:@11380.4]
  assign _T_29255 = _T_29254 | _T_29224; // @[Mux.scala 19:72:@11381.4]
  assign _T_29256 = _T_29255 | _T_29233; // @[Mux.scala 19:72:@11382.4]
  assign _T_29257 = _T_29256 | _T_29242; // @[Mux.scala 19:72:@11383.4]
  assign _T_29258 = _T_29257 | _T_29251; // @[Mux.scala 19:72:@11384.4]
  assign outputPriorityPorts_2_0 = _T_29258[0]; // @[Mux.scala 19:72:@11388.4]
  assign outputPriorityPorts_2_1 = _T_29258[1]; // @[Mux.scala 19:72:@11390.4]
  assign outputPriorityPorts_2_2 = _T_29258[2]; // @[Mux.scala 19:72:@11392.4]
  assign outputPriorityPorts_2_3 = _T_29258[3]; // @[Mux.scala 19:72:@11394.4]
  assign outputPriorityPorts_2_4 = _T_29258[4]; // @[Mux.scala 19:72:@11396.4]
  assign outputPriorityPorts_2_5 = _T_29258[5]; // @[Mux.scala 19:72:@11398.4]
  assign outputPriorityPorts_2_6 = _T_29258[6]; // @[Mux.scala 19:72:@11400.4]
  assign outputPriorityPorts_2_7 = _T_29258[7]; // @[Mux.scala 19:72:@11402.4]
  assign _T_29338 = entriesPorts_3_0 & _T_26091; // @[LoadQueue.scala 298:83:@11413.4]
  assign _T_29341 = entriesPorts_3_1 & _T_26094; // @[LoadQueue.scala 298:83:@11415.4]
  assign _T_29344 = entriesPorts_3_2 & _T_26097; // @[LoadQueue.scala 298:83:@11417.4]
  assign _T_29347 = entriesPorts_3_3 & _T_26100; // @[LoadQueue.scala 298:83:@11419.4]
  assign _T_29350 = entriesPorts_3_4 & _T_26103; // @[LoadQueue.scala 298:83:@11421.4]
  assign _T_29353 = entriesPorts_3_5 & _T_26106; // @[LoadQueue.scala 298:83:@11423.4]
  assign _T_29356 = entriesPorts_3_6 & _T_26109; // @[LoadQueue.scala 298:83:@11425.4]
  assign _T_29359 = entriesPorts_3_7 & _T_26112; // @[LoadQueue.scala 298:83:@11427.4]
  assign _T_29410 = _T_29359 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11457.4]
  assign _T_29411 = _T_29356 ? 8'h40 : _T_29410; // @[Mux.scala 31:69:@11458.4]
  assign _T_29412 = _T_29353 ? 8'h20 : _T_29411; // @[Mux.scala 31:69:@11459.4]
  assign _T_29413 = _T_29350 ? 8'h10 : _T_29412; // @[Mux.scala 31:69:@11460.4]
  assign _T_29414 = _T_29347 ? 8'h8 : _T_29413; // @[Mux.scala 31:69:@11461.4]
  assign _T_29415 = _T_29344 ? 8'h4 : _T_29414; // @[Mux.scala 31:69:@11462.4]
  assign _T_29416 = _T_29341 ? 8'h2 : _T_29415; // @[Mux.scala 31:69:@11463.4]
  assign _T_29417 = _T_29338 ? 8'h1 : _T_29416; // @[Mux.scala 31:69:@11464.4]
  assign _T_29418 = _T_29417[0]; // @[OneHot.scala 66:30:@11465.4]
  assign _T_29419 = _T_29417[1]; // @[OneHot.scala 66:30:@11466.4]
  assign _T_29420 = _T_29417[2]; // @[OneHot.scala 66:30:@11467.4]
  assign _T_29421 = _T_29417[3]; // @[OneHot.scala 66:30:@11468.4]
  assign _T_29422 = _T_29417[4]; // @[OneHot.scala 66:30:@11469.4]
  assign _T_29423 = _T_29417[5]; // @[OneHot.scala 66:30:@11470.4]
  assign _T_29424 = _T_29417[6]; // @[OneHot.scala 66:30:@11471.4]
  assign _T_29425 = _T_29417[7]; // @[OneHot.scala 66:30:@11472.4]
  assign _T_29450 = _T_29338 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11482.4]
  assign _T_29451 = _T_29359 ? 8'h40 : _T_29450; // @[Mux.scala 31:69:@11483.4]
  assign _T_29452 = _T_29356 ? 8'h20 : _T_29451; // @[Mux.scala 31:69:@11484.4]
  assign _T_29453 = _T_29353 ? 8'h10 : _T_29452; // @[Mux.scala 31:69:@11485.4]
  assign _T_29454 = _T_29350 ? 8'h8 : _T_29453; // @[Mux.scala 31:69:@11486.4]
  assign _T_29455 = _T_29347 ? 8'h4 : _T_29454; // @[Mux.scala 31:69:@11487.4]
  assign _T_29456 = _T_29344 ? 8'h2 : _T_29455; // @[Mux.scala 31:69:@11488.4]
  assign _T_29457 = _T_29341 ? 8'h1 : _T_29456; // @[Mux.scala 31:69:@11489.4]
  assign _T_29458 = _T_29457[0]; // @[OneHot.scala 66:30:@11490.4]
  assign _T_29459 = _T_29457[1]; // @[OneHot.scala 66:30:@11491.4]
  assign _T_29460 = _T_29457[2]; // @[OneHot.scala 66:30:@11492.4]
  assign _T_29461 = _T_29457[3]; // @[OneHot.scala 66:30:@11493.4]
  assign _T_29462 = _T_29457[4]; // @[OneHot.scala 66:30:@11494.4]
  assign _T_29463 = _T_29457[5]; // @[OneHot.scala 66:30:@11495.4]
  assign _T_29464 = _T_29457[6]; // @[OneHot.scala 66:30:@11496.4]
  assign _T_29465 = _T_29457[7]; // @[OneHot.scala 66:30:@11497.4]
  assign _T_29490 = _T_29341 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11507.4]
  assign _T_29491 = _T_29338 ? 8'h40 : _T_29490; // @[Mux.scala 31:69:@11508.4]
  assign _T_29492 = _T_29359 ? 8'h20 : _T_29491; // @[Mux.scala 31:69:@11509.4]
  assign _T_29493 = _T_29356 ? 8'h10 : _T_29492; // @[Mux.scala 31:69:@11510.4]
  assign _T_29494 = _T_29353 ? 8'h8 : _T_29493; // @[Mux.scala 31:69:@11511.4]
  assign _T_29495 = _T_29350 ? 8'h4 : _T_29494; // @[Mux.scala 31:69:@11512.4]
  assign _T_29496 = _T_29347 ? 8'h2 : _T_29495; // @[Mux.scala 31:69:@11513.4]
  assign _T_29497 = _T_29344 ? 8'h1 : _T_29496; // @[Mux.scala 31:69:@11514.4]
  assign _T_29498 = _T_29497[0]; // @[OneHot.scala 66:30:@11515.4]
  assign _T_29499 = _T_29497[1]; // @[OneHot.scala 66:30:@11516.4]
  assign _T_29500 = _T_29497[2]; // @[OneHot.scala 66:30:@11517.4]
  assign _T_29501 = _T_29497[3]; // @[OneHot.scala 66:30:@11518.4]
  assign _T_29502 = _T_29497[4]; // @[OneHot.scala 66:30:@11519.4]
  assign _T_29503 = _T_29497[5]; // @[OneHot.scala 66:30:@11520.4]
  assign _T_29504 = _T_29497[6]; // @[OneHot.scala 66:30:@11521.4]
  assign _T_29505 = _T_29497[7]; // @[OneHot.scala 66:30:@11522.4]
  assign _T_29530 = _T_29344 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11532.4]
  assign _T_29531 = _T_29341 ? 8'h40 : _T_29530; // @[Mux.scala 31:69:@11533.4]
  assign _T_29532 = _T_29338 ? 8'h20 : _T_29531; // @[Mux.scala 31:69:@11534.4]
  assign _T_29533 = _T_29359 ? 8'h10 : _T_29532; // @[Mux.scala 31:69:@11535.4]
  assign _T_29534 = _T_29356 ? 8'h8 : _T_29533; // @[Mux.scala 31:69:@11536.4]
  assign _T_29535 = _T_29353 ? 8'h4 : _T_29534; // @[Mux.scala 31:69:@11537.4]
  assign _T_29536 = _T_29350 ? 8'h2 : _T_29535; // @[Mux.scala 31:69:@11538.4]
  assign _T_29537 = _T_29347 ? 8'h1 : _T_29536; // @[Mux.scala 31:69:@11539.4]
  assign _T_29538 = _T_29537[0]; // @[OneHot.scala 66:30:@11540.4]
  assign _T_29539 = _T_29537[1]; // @[OneHot.scala 66:30:@11541.4]
  assign _T_29540 = _T_29537[2]; // @[OneHot.scala 66:30:@11542.4]
  assign _T_29541 = _T_29537[3]; // @[OneHot.scala 66:30:@11543.4]
  assign _T_29542 = _T_29537[4]; // @[OneHot.scala 66:30:@11544.4]
  assign _T_29543 = _T_29537[5]; // @[OneHot.scala 66:30:@11545.4]
  assign _T_29544 = _T_29537[6]; // @[OneHot.scala 66:30:@11546.4]
  assign _T_29545 = _T_29537[7]; // @[OneHot.scala 66:30:@11547.4]
  assign _T_29570 = _T_29347 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11557.4]
  assign _T_29571 = _T_29344 ? 8'h40 : _T_29570; // @[Mux.scala 31:69:@11558.4]
  assign _T_29572 = _T_29341 ? 8'h20 : _T_29571; // @[Mux.scala 31:69:@11559.4]
  assign _T_29573 = _T_29338 ? 8'h10 : _T_29572; // @[Mux.scala 31:69:@11560.4]
  assign _T_29574 = _T_29359 ? 8'h8 : _T_29573; // @[Mux.scala 31:69:@11561.4]
  assign _T_29575 = _T_29356 ? 8'h4 : _T_29574; // @[Mux.scala 31:69:@11562.4]
  assign _T_29576 = _T_29353 ? 8'h2 : _T_29575; // @[Mux.scala 31:69:@11563.4]
  assign _T_29577 = _T_29350 ? 8'h1 : _T_29576; // @[Mux.scala 31:69:@11564.4]
  assign _T_29578 = _T_29577[0]; // @[OneHot.scala 66:30:@11565.4]
  assign _T_29579 = _T_29577[1]; // @[OneHot.scala 66:30:@11566.4]
  assign _T_29580 = _T_29577[2]; // @[OneHot.scala 66:30:@11567.4]
  assign _T_29581 = _T_29577[3]; // @[OneHot.scala 66:30:@11568.4]
  assign _T_29582 = _T_29577[4]; // @[OneHot.scala 66:30:@11569.4]
  assign _T_29583 = _T_29577[5]; // @[OneHot.scala 66:30:@11570.4]
  assign _T_29584 = _T_29577[6]; // @[OneHot.scala 66:30:@11571.4]
  assign _T_29585 = _T_29577[7]; // @[OneHot.scala 66:30:@11572.4]
  assign _T_29610 = _T_29350 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11582.4]
  assign _T_29611 = _T_29347 ? 8'h40 : _T_29610; // @[Mux.scala 31:69:@11583.4]
  assign _T_29612 = _T_29344 ? 8'h20 : _T_29611; // @[Mux.scala 31:69:@11584.4]
  assign _T_29613 = _T_29341 ? 8'h10 : _T_29612; // @[Mux.scala 31:69:@11585.4]
  assign _T_29614 = _T_29338 ? 8'h8 : _T_29613; // @[Mux.scala 31:69:@11586.4]
  assign _T_29615 = _T_29359 ? 8'h4 : _T_29614; // @[Mux.scala 31:69:@11587.4]
  assign _T_29616 = _T_29356 ? 8'h2 : _T_29615; // @[Mux.scala 31:69:@11588.4]
  assign _T_29617 = _T_29353 ? 8'h1 : _T_29616; // @[Mux.scala 31:69:@11589.4]
  assign _T_29618 = _T_29617[0]; // @[OneHot.scala 66:30:@11590.4]
  assign _T_29619 = _T_29617[1]; // @[OneHot.scala 66:30:@11591.4]
  assign _T_29620 = _T_29617[2]; // @[OneHot.scala 66:30:@11592.4]
  assign _T_29621 = _T_29617[3]; // @[OneHot.scala 66:30:@11593.4]
  assign _T_29622 = _T_29617[4]; // @[OneHot.scala 66:30:@11594.4]
  assign _T_29623 = _T_29617[5]; // @[OneHot.scala 66:30:@11595.4]
  assign _T_29624 = _T_29617[6]; // @[OneHot.scala 66:30:@11596.4]
  assign _T_29625 = _T_29617[7]; // @[OneHot.scala 66:30:@11597.4]
  assign _T_29650 = _T_29353 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11607.4]
  assign _T_29651 = _T_29350 ? 8'h40 : _T_29650; // @[Mux.scala 31:69:@11608.4]
  assign _T_29652 = _T_29347 ? 8'h20 : _T_29651; // @[Mux.scala 31:69:@11609.4]
  assign _T_29653 = _T_29344 ? 8'h10 : _T_29652; // @[Mux.scala 31:69:@11610.4]
  assign _T_29654 = _T_29341 ? 8'h8 : _T_29653; // @[Mux.scala 31:69:@11611.4]
  assign _T_29655 = _T_29338 ? 8'h4 : _T_29654; // @[Mux.scala 31:69:@11612.4]
  assign _T_29656 = _T_29359 ? 8'h2 : _T_29655; // @[Mux.scala 31:69:@11613.4]
  assign _T_29657 = _T_29356 ? 8'h1 : _T_29656; // @[Mux.scala 31:69:@11614.4]
  assign _T_29658 = _T_29657[0]; // @[OneHot.scala 66:30:@11615.4]
  assign _T_29659 = _T_29657[1]; // @[OneHot.scala 66:30:@11616.4]
  assign _T_29660 = _T_29657[2]; // @[OneHot.scala 66:30:@11617.4]
  assign _T_29661 = _T_29657[3]; // @[OneHot.scala 66:30:@11618.4]
  assign _T_29662 = _T_29657[4]; // @[OneHot.scala 66:30:@11619.4]
  assign _T_29663 = _T_29657[5]; // @[OneHot.scala 66:30:@11620.4]
  assign _T_29664 = _T_29657[6]; // @[OneHot.scala 66:30:@11621.4]
  assign _T_29665 = _T_29657[7]; // @[OneHot.scala 66:30:@11622.4]
  assign _T_29690 = _T_29356 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11632.4]
  assign _T_29691 = _T_29353 ? 8'h40 : _T_29690; // @[Mux.scala 31:69:@11633.4]
  assign _T_29692 = _T_29350 ? 8'h20 : _T_29691; // @[Mux.scala 31:69:@11634.4]
  assign _T_29693 = _T_29347 ? 8'h10 : _T_29692; // @[Mux.scala 31:69:@11635.4]
  assign _T_29694 = _T_29344 ? 8'h8 : _T_29693; // @[Mux.scala 31:69:@11636.4]
  assign _T_29695 = _T_29341 ? 8'h4 : _T_29694; // @[Mux.scala 31:69:@11637.4]
  assign _T_29696 = _T_29338 ? 8'h2 : _T_29695; // @[Mux.scala 31:69:@11638.4]
  assign _T_29697 = _T_29359 ? 8'h1 : _T_29696; // @[Mux.scala 31:69:@11639.4]
  assign _T_29698 = _T_29697[0]; // @[OneHot.scala 66:30:@11640.4]
  assign _T_29699 = _T_29697[1]; // @[OneHot.scala 66:30:@11641.4]
  assign _T_29700 = _T_29697[2]; // @[OneHot.scala 66:30:@11642.4]
  assign _T_29701 = _T_29697[3]; // @[OneHot.scala 66:30:@11643.4]
  assign _T_29702 = _T_29697[4]; // @[OneHot.scala 66:30:@11644.4]
  assign _T_29703 = _T_29697[5]; // @[OneHot.scala 66:30:@11645.4]
  assign _T_29704 = _T_29697[6]; // @[OneHot.scala 66:30:@11646.4]
  assign _T_29705 = _T_29697[7]; // @[OneHot.scala 66:30:@11647.4]
  assign _T_29746 = {_T_29425,_T_29424,_T_29423,_T_29422,_T_29421,_T_29420,_T_29419,_T_29418}; // @[Mux.scala 19:72:@11663.4]
  assign _T_29748 = _T_24176 ? _T_29746 : 8'h0; // @[Mux.scala 19:72:@11664.4]
  assign _T_29755 = {_T_29464,_T_29463,_T_29462,_T_29461,_T_29460,_T_29459,_T_29458,_T_29465}; // @[Mux.scala 19:72:@11671.4]
  assign _T_29757 = _T_24177 ? _T_29755 : 8'h0; // @[Mux.scala 19:72:@11672.4]
  assign _T_29764 = {_T_29503,_T_29502,_T_29501,_T_29500,_T_29499,_T_29498,_T_29505,_T_29504}; // @[Mux.scala 19:72:@11679.4]
  assign _T_29766 = _T_24178 ? _T_29764 : 8'h0; // @[Mux.scala 19:72:@11680.4]
  assign _T_29773 = {_T_29542,_T_29541,_T_29540,_T_29539,_T_29538,_T_29545,_T_29544,_T_29543}; // @[Mux.scala 19:72:@11687.4]
  assign _T_29775 = _T_24179 ? _T_29773 : 8'h0; // @[Mux.scala 19:72:@11688.4]
  assign _T_29782 = {_T_29581,_T_29580,_T_29579,_T_29578,_T_29585,_T_29584,_T_29583,_T_29582}; // @[Mux.scala 19:72:@11695.4]
  assign _T_29784 = _T_24180 ? _T_29782 : 8'h0; // @[Mux.scala 19:72:@11696.4]
  assign _T_29791 = {_T_29620,_T_29619,_T_29618,_T_29625,_T_29624,_T_29623,_T_29622,_T_29621}; // @[Mux.scala 19:72:@11703.4]
  assign _T_29793 = _T_24181 ? _T_29791 : 8'h0; // @[Mux.scala 19:72:@11704.4]
  assign _T_29800 = {_T_29659,_T_29658,_T_29665,_T_29664,_T_29663,_T_29662,_T_29661,_T_29660}; // @[Mux.scala 19:72:@11711.4]
  assign _T_29802 = _T_24182 ? _T_29800 : 8'h0; // @[Mux.scala 19:72:@11712.4]
  assign _T_29809 = {_T_29698,_T_29705,_T_29704,_T_29703,_T_29702,_T_29701,_T_29700,_T_29699}; // @[Mux.scala 19:72:@11719.4]
  assign _T_29811 = _T_24183 ? _T_29809 : 8'h0; // @[Mux.scala 19:72:@11720.4]
  assign _T_29812 = _T_29748 | _T_29757; // @[Mux.scala 19:72:@11721.4]
  assign _T_29813 = _T_29812 | _T_29766; // @[Mux.scala 19:72:@11722.4]
  assign _T_29814 = _T_29813 | _T_29775; // @[Mux.scala 19:72:@11723.4]
  assign _T_29815 = _T_29814 | _T_29784; // @[Mux.scala 19:72:@11724.4]
  assign _T_29816 = _T_29815 | _T_29793; // @[Mux.scala 19:72:@11725.4]
  assign _T_29817 = _T_29816 | _T_29802; // @[Mux.scala 19:72:@11726.4]
  assign _T_29818 = _T_29817 | _T_29811; // @[Mux.scala 19:72:@11727.4]
  assign inputPriorityPorts_3_0 = _T_29818[0]; // @[Mux.scala 19:72:@11731.4]
  assign inputPriorityPorts_3_1 = _T_29818[1]; // @[Mux.scala 19:72:@11733.4]
  assign inputPriorityPorts_3_2 = _T_29818[2]; // @[Mux.scala 19:72:@11735.4]
  assign inputPriorityPorts_3_3 = _T_29818[3]; // @[Mux.scala 19:72:@11737.4]
  assign inputPriorityPorts_3_4 = _T_29818[4]; // @[Mux.scala 19:72:@11739.4]
  assign inputPriorityPorts_3_5 = _T_29818[5]; // @[Mux.scala 19:72:@11741.4]
  assign inputPriorityPorts_3_6 = _T_29818[6]; // @[Mux.scala 19:72:@11743.4]
  assign inputPriorityPorts_3_7 = _T_29818[7]; // @[Mux.scala 19:72:@11745.4]
  assign _T_29932 = entriesPorts_3_7 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11775.4]
  assign _T_29933 = entriesPorts_3_6 ? 8'h40 : _T_29932; // @[Mux.scala 31:69:@11776.4]
  assign _T_29934 = entriesPorts_3_5 ? 8'h20 : _T_29933; // @[Mux.scala 31:69:@11777.4]
  assign _T_29935 = entriesPorts_3_4 ? 8'h10 : _T_29934; // @[Mux.scala 31:69:@11778.4]
  assign _T_29936 = entriesPorts_3_3 ? 8'h8 : _T_29935; // @[Mux.scala 31:69:@11779.4]
  assign _T_29937 = entriesPorts_3_2 ? 8'h4 : _T_29936; // @[Mux.scala 31:69:@11780.4]
  assign _T_29938 = entriesPorts_3_1 ? 8'h2 : _T_29937; // @[Mux.scala 31:69:@11781.4]
  assign _T_29939 = entriesPorts_3_0 ? 8'h1 : _T_29938; // @[Mux.scala 31:69:@11782.4]
  assign _T_29940 = _T_29939[0]; // @[OneHot.scala 66:30:@11783.4]
  assign _T_29941 = _T_29939[1]; // @[OneHot.scala 66:30:@11784.4]
  assign _T_29942 = _T_29939[2]; // @[OneHot.scala 66:30:@11785.4]
  assign _T_29943 = _T_29939[3]; // @[OneHot.scala 66:30:@11786.4]
  assign _T_29944 = _T_29939[4]; // @[OneHot.scala 66:30:@11787.4]
  assign _T_29945 = _T_29939[5]; // @[OneHot.scala 66:30:@11788.4]
  assign _T_29946 = _T_29939[6]; // @[OneHot.scala 66:30:@11789.4]
  assign _T_29947 = _T_29939[7]; // @[OneHot.scala 66:30:@11790.4]
  assign _T_29972 = entriesPorts_3_0 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11800.4]
  assign _T_29973 = entriesPorts_3_7 ? 8'h40 : _T_29972; // @[Mux.scala 31:69:@11801.4]
  assign _T_29974 = entriesPorts_3_6 ? 8'h20 : _T_29973; // @[Mux.scala 31:69:@11802.4]
  assign _T_29975 = entriesPorts_3_5 ? 8'h10 : _T_29974; // @[Mux.scala 31:69:@11803.4]
  assign _T_29976 = entriesPorts_3_4 ? 8'h8 : _T_29975; // @[Mux.scala 31:69:@11804.4]
  assign _T_29977 = entriesPorts_3_3 ? 8'h4 : _T_29976; // @[Mux.scala 31:69:@11805.4]
  assign _T_29978 = entriesPorts_3_2 ? 8'h2 : _T_29977; // @[Mux.scala 31:69:@11806.4]
  assign _T_29979 = entriesPorts_3_1 ? 8'h1 : _T_29978; // @[Mux.scala 31:69:@11807.4]
  assign _T_29980 = _T_29979[0]; // @[OneHot.scala 66:30:@11808.4]
  assign _T_29981 = _T_29979[1]; // @[OneHot.scala 66:30:@11809.4]
  assign _T_29982 = _T_29979[2]; // @[OneHot.scala 66:30:@11810.4]
  assign _T_29983 = _T_29979[3]; // @[OneHot.scala 66:30:@11811.4]
  assign _T_29984 = _T_29979[4]; // @[OneHot.scala 66:30:@11812.4]
  assign _T_29985 = _T_29979[5]; // @[OneHot.scala 66:30:@11813.4]
  assign _T_29986 = _T_29979[6]; // @[OneHot.scala 66:30:@11814.4]
  assign _T_29987 = _T_29979[7]; // @[OneHot.scala 66:30:@11815.4]
  assign _T_30012 = entriesPorts_3_1 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11825.4]
  assign _T_30013 = entriesPorts_3_0 ? 8'h40 : _T_30012; // @[Mux.scala 31:69:@11826.4]
  assign _T_30014 = entriesPorts_3_7 ? 8'h20 : _T_30013; // @[Mux.scala 31:69:@11827.4]
  assign _T_30015 = entriesPorts_3_6 ? 8'h10 : _T_30014; // @[Mux.scala 31:69:@11828.4]
  assign _T_30016 = entriesPorts_3_5 ? 8'h8 : _T_30015; // @[Mux.scala 31:69:@11829.4]
  assign _T_30017 = entriesPorts_3_4 ? 8'h4 : _T_30016; // @[Mux.scala 31:69:@11830.4]
  assign _T_30018 = entriesPorts_3_3 ? 8'h2 : _T_30017; // @[Mux.scala 31:69:@11831.4]
  assign _T_30019 = entriesPorts_3_2 ? 8'h1 : _T_30018; // @[Mux.scala 31:69:@11832.4]
  assign _T_30020 = _T_30019[0]; // @[OneHot.scala 66:30:@11833.4]
  assign _T_30021 = _T_30019[1]; // @[OneHot.scala 66:30:@11834.4]
  assign _T_30022 = _T_30019[2]; // @[OneHot.scala 66:30:@11835.4]
  assign _T_30023 = _T_30019[3]; // @[OneHot.scala 66:30:@11836.4]
  assign _T_30024 = _T_30019[4]; // @[OneHot.scala 66:30:@11837.4]
  assign _T_30025 = _T_30019[5]; // @[OneHot.scala 66:30:@11838.4]
  assign _T_30026 = _T_30019[6]; // @[OneHot.scala 66:30:@11839.4]
  assign _T_30027 = _T_30019[7]; // @[OneHot.scala 66:30:@11840.4]
  assign _T_30052 = entriesPorts_3_2 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11850.4]
  assign _T_30053 = entriesPorts_3_1 ? 8'h40 : _T_30052; // @[Mux.scala 31:69:@11851.4]
  assign _T_30054 = entriesPorts_3_0 ? 8'h20 : _T_30053; // @[Mux.scala 31:69:@11852.4]
  assign _T_30055 = entriesPorts_3_7 ? 8'h10 : _T_30054; // @[Mux.scala 31:69:@11853.4]
  assign _T_30056 = entriesPorts_3_6 ? 8'h8 : _T_30055; // @[Mux.scala 31:69:@11854.4]
  assign _T_30057 = entriesPorts_3_5 ? 8'h4 : _T_30056; // @[Mux.scala 31:69:@11855.4]
  assign _T_30058 = entriesPorts_3_4 ? 8'h2 : _T_30057; // @[Mux.scala 31:69:@11856.4]
  assign _T_30059 = entriesPorts_3_3 ? 8'h1 : _T_30058; // @[Mux.scala 31:69:@11857.4]
  assign _T_30060 = _T_30059[0]; // @[OneHot.scala 66:30:@11858.4]
  assign _T_30061 = _T_30059[1]; // @[OneHot.scala 66:30:@11859.4]
  assign _T_30062 = _T_30059[2]; // @[OneHot.scala 66:30:@11860.4]
  assign _T_30063 = _T_30059[3]; // @[OneHot.scala 66:30:@11861.4]
  assign _T_30064 = _T_30059[4]; // @[OneHot.scala 66:30:@11862.4]
  assign _T_30065 = _T_30059[5]; // @[OneHot.scala 66:30:@11863.4]
  assign _T_30066 = _T_30059[6]; // @[OneHot.scala 66:30:@11864.4]
  assign _T_30067 = _T_30059[7]; // @[OneHot.scala 66:30:@11865.4]
  assign _T_30092 = entriesPorts_3_3 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11875.4]
  assign _T_30093 = entriesPorts_3_2 ? 8'h40 : _T_30092; // @[Mux.scala 31:69:@11876.4]
  assign _T_30094 = entriesPorts_3_1 ? 8'h20 : _T_30093; // @[Mux.scala 31:69:@11877.4]
  assign _T_30095 = entriesPorts_3_0 ? 8'h10 : _T_30094; // @[Mux.scala 31:69:@11878.4]
  assign _T_30096 = entriesPorts_3_7 ? 8'h8 : _T_30095; // @[Mux.scala 31:69:@11879.4]
  assign _T_30097 = entriesPorts_3_6 ? 8'h4 : _T_30096; // @[Mux.scala 31:69:@11880.4]
  assign _T_30098 = entriesPorts_3_5 ? 8'h2 : _T_30097; // @[Mux.scala 31:69:@11881.4]
  assign _T_30099 = entriesPorts_3_4 ? 8'h1 : _T_30098; // @[Mux.scala 31:69:@11882.4]
  assign _T_30100 = _T_30099[0]; // @[OneHot.scala 66:30:@11883.4]
  assign _T_30101 = _T_30099[1]; // @[OneHot.scala 66:30:@11884.4]
  assign _T_30102 = _T_30099[2]; // @[OneHot.scala 66:30:@11885.4]
  assign _T_30103 = _T_30099[3]; // @[OneHot.scala 66:30:@11886.4]
  assign _T_30104 = _T_30099[4]; // @[OneHot.scala 66:30:@11887.4]
  assign _T_30105 = _T_30099[5]; // @[OneHot.scala 66:30:@11888.4]
  assign _T_30106 = _T_30099[6]; // @[OneHot.scala 66:30:@11889.4]
  assign _T_30107 = _T_30099[7]; // @[OneHot.scala 66:30:@11890.4]
  assign _T_30132 = entriesPorts_3_4 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11900.4]
  assign _T_30133 = entriesPorts_3_3 ? 8'h40 : _T_30132; // @[Mux.scala 31:69:@11901.4]
  assign _T_30134 = entriesPorts_3_2 ? 8'h20 : _T_30133; // @[Mux.scala 31:69:@11902.4]
  assign _T_30135 = entriesPorts_3_1 ? 8'h10 : _T_30134; // @[Mux.scala 31:69:@11903.4]
  assign _T_30136 = entriesPorts_3_0 ? 8'h8 : _T_30135; // @[Mux.scala 31:69:@11904.4]
  assign _T_30137 = entriesPorts_3_7 ? 8'h4 : _T_30136; // @[Mux.scala 31:69:@11905.4]
  assign _T_30138 = entriesPorts_3_6 ? 8'h2 : _T_30137; // @[Mux.scala 31:69:@11906.4]
  assign _T_30139 = entriesPorts_3_5 ? 8'h1 : _T_30138; // @[Mux.scala 31:69:@11907.4]
  assign _T_30140 = _T_30139[0]; // @[OneHot.scala 66:30:@11908.4]
  assign _T_30141 = _T_30139[1]; // @[OneHot.scala 66:30:@11909.4]
  assign _T_30142 = _T_30139[2]; // @[OneHot.scala 66:30:@11910.4]
  assign _T_30143 = _T_30139[3]; // @[OneHot.scala 66:30:@11911.4]
  assign _T_30144 = _T_30139[4]; // @[OneHot.scala 66:30:@11912.4]
  assign _T_30145 = _T_30139[5]; // @[OneHot.scala 66:30:@11913.4]
  assign _T_30146 = _T_30139[6]; // @[OneHot.scala 66:30:@11914.4]
  assign _T_30147 = _T_30139[7]; // @[OneHot.scala 66:30:@11915.4]
  assign _T_30172 = entriesPorts_3_5 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11925.4]
  assign _T_30173 = entriesPorts_3_4 ? 8'h40 : _T_30172; // @[Mux.scala 31:69:@11926.4]
  assign _T_30174 = entriesPorts_3_3 ? 8'h20 : _T_30173; // @[Mux.scala 31:69:@11927.4]
  assign _T_30175 = entriesPorts_3_2 ? 8'h10 : _T_30174; // @[Mux.scala 31:69:@11928.4]
  assign _T_30176 = entriesPorts_3_1 ? 8'h8 : _T_30175; // @[Mux.scala 31:69:@11929.4]
  assign _T_30177 = entriesPorts_3_0 ? 8'h4 : _T_30176; // @[Mux.scala 31:69:@11930.4]
  assign _T_30178 = entriesPorts_3_7 ? 8'h2 : _T_30177; // @[Mux.scala 31:69:@11931.4]
  assign _T_30179 = entriesPorts_3_6 ? 8'h1 : _T_30178; // @[Mux.scala 31:69:@11932.4]
  assign _T_30180 = _T_30179[0]; // @[OneHot.scala 66:30:@11933.4]
  assign _T_30181 = _T_30179[1]; // @[OneHot.scala 66:30:@11934.4]
  assign _T_30182 = _T_30179[2]; // @[OneHot.scala 66:30:@11935.4]
  assign _T_30183 = _T_30179[3]; // @[OneHot.scala 66:30:@11936.4]
  assign _T_30184 = _T_30179[4]; // @[OneHot.scala 66:30:@11937.4]
  assign _T_30185 = _T_30179[5]; // @[OneHot.scala 66:30:@11938.4]
  assign _T_30186 = _T_30179[6]; // @[OneHot.scala 66:30:@11939.4]
  assign _T_30187 = _T_30179[7]; // @[OneHot.scala 66:30:@11940.4]
  assign _T_30212 = entriesPorts_3_6 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11950.4]
  assign _T_30213 = entriesPorts_3_5 ? 8'h40 : _T_30212; // @[Mux.scala 31:69:@11951.4]
  assign _T_30214 = entriesPorts_3_4 ? 8'h20 : _T_30213; // @[Mux.scala 31:69:@11952.4]
  assign _T_30215 = entriesPorts_3_3 ? 8'h10 : _T_30214; // @[Mux.scala 31:69:@11953.4]
  assign _T_30216 = entriesPorts_3_2 ? 8'h8 : _T_30215; // @[Mux.scala 31:69:@11954.4]
  assign _T_30217 = entriesPorts_3_1 ? 8'h4 : _T_30216; // @[Mux.scala 31:69:@11955.4]
  assign _T_30218 = entriesPorts_3_0 ? 8'h2 : _T_30217; // @[Mux.scala 31:69:@11956.4]
  assign _T_30219 = entriesPorts_3_7 ? 8'h1 : _T_30218; // @[Mux.scala 31:69:@11957.4]
  assign _T_30220 = _T_30219[0]; // @[OneHot.scala 66:30:@11958.4]
  assign _T_30221 = _T_30219[1]; // @[OneHot.scala 66:30:@11959.4]
  assign _T_30222 = _T_30219[2]; // @[OneHot.scala 66:30:@11960.4]
  assign _T_30223 = _T_30219[3]; // @[OneHot.scala 66:30:@11961.4]
  assign _T_30224 = _T_30219[4]; // @[OneHot.scala 66:30:@11962.4]
  assign _T_30225 = _T_30219[5]; // @[OneHot.scala 66:30:@11963.4]
  assign _T_30226 = _T_30219[6]; // @[OneHot.scala 66:30:@11964.4]
  assign _T_30227 = _T_30219[7]; // @[OneHot.scala 66:30:@11965.4]
  assign _T_30268 = {_T_29947,_T_29946,_T_29945,_T_29944,_T_29943,_T_29942,_T_29941,_T_29940}; // @[Mux.scala 19:72:@11981.4]
  assign _T_30270 = _T_24176 ? _T_30268 : 8'h0; // @[Mux.scala 19:72:@11982.4]
  assign _T_30277 = {_T_29986,_T_29985,_T_29984,_T_29983,_T_29982,_T_29981,_T_29980,_T_29987}; // @[Mux.scala 19:72:@11989.4]
  assign _T_30279 = _T_24177 ? _T_30277 : 8'h0; // @[Mux.scala 19:72:@11990.4]
  assign _T_30286 = {_T_30025,_T_30024,_T_30023,_T_30022,_T_30021,_T_30020,_T_30027,_T_30026}; // @[Mux.scala 19:72:@11997.4]
  assign _T_30288 = _T_24178 ? _T_30286 : 8'h0; // @[Mux.scala 19:72:@11998.4]
  assign _T_30295 = {_T_30064,_T_30063,_T_30062,_T_30061,_T_30060,_T_30067,_T_30066,_T_30065}; // @[Mux.scala 19:72:@12005.4]
  assign _T_30297 = _T_24179 ? _T_30295 : 8'h0; // @[Mux.scala 19:72:@12006.4]
  assign _T_30304 = {_T_30103,_T_30102,_T_30101,_T_30100,_T_30107,_T_30106,_T_30105,_T_30104}; // @[Mux.scala 19:72:@12013.4]
  assign _T_30306 = _T_24180 ? _T_30304 : 8'h0; // @[Mux.scala 19:72:@12014.4]
  assign _T_30313 = {_T_30142,_T_30141,_T_30140,_T_30147,_T_30146,_T_30145,_T_30144,_T_30143}; // @[Mux.scala 19:72:@12021.4]
  assign _T_30315 = _T_24181 ? _T_30313 : 8'h0; // @[Mux.scala 19:72:@12022.4]
  assign _T_30322 = {_T_30181,_T_30180,_T_30187,_T_30186,_T_30185,_T_30184,_T_30183,_T_30182}; // @[Mux.scala 19:72:@12029.4]
  assign _T_30324 = _T_24182 ? _T_30322 : 8'h0; // @[Mux.scala 19:72:@12030.4]
  assign _T_30331 = {_T_30220,_T_30227,_T_30226,_T_30225,_T_30224,_T_30223,_T_30222,_T_30221}; // @[Mux.scala 19:72:@12037.4]
  assign _T_30333 = _T_24183 ? _T_30331 : 8'h0; // @[Mux.scala 19:72:@12038.4]
  assign _T_30334 = _T_30270 | _T_30279; // @[Mux.scala 19:72:@12039.4]
  assign _T_30335 = _T_30334 | _T_30288; // @[Mux.scala 19:72:@12040.4]
  assign _T_30336 = _T_30335 | _T_30297; // @[Mux.scala 19:72:@12041.4]
  assign _T_30337 = _T_30336 | _T_30306; // @[Mux.scala 19:72:@12042.4]
  assign _T_30338 = _T_30337 | _T_30315; // @[Mux.scala 19:72:@12043.4]
  assign _T_30339 = _T_30338 | _T_30324; // @[Mux.scala 19:72:@12044.4]
  assign _T_30340 = _T_30339 | _T_30333; // @[Mux.scala 19:72:@12045.4]
  assign outputPriorityPorts_3_0 = _T_30340[0]; // @[Mux.scala 19:72:@12049.4]
  assign outputPriorityPorts_3_1 = _T_30340[1]; // @[Mux.scala 19:72:@12051.4]
  assign outputPriorityPorts_3_2 = _T_30340[2]; // @[Mux.scala 19:72:@12053.4]
  assign outputPriorityPorts_3_3 = _T_30340[3]; // @[Mux.scala 19:72:@12055.4]
  assign outputPriorityPorts_3_4 = _T_30340[4]; // @[Mux.scala 19:72:@12057.4]
  assign outputPriorityPorts_3_5 = _T_30340[5]; // @[Mux.scala 19:72:@12059.4]
  assign outputPriorityPorts_3_6 = _T_30340[6]; // @[Mux.scala 19:72:@12061.4]
  assign outputPriorityPorts_3_7 = _T_30340[7]; // @[Mux.scala 19:72:@12063.4]
  assign _T_30420 = entriesPorts_4_0 & _T_26091; // @[LoadQueue.scala 298:83:@12074.4]
  assign _T_30423 = entriesPorts_4_1 & _T_26094; // @[LoadQueue.scala 298:83:@12076.4]
  assign _T_30426 = entriesPorts_4_2 & _T_26097; // @[LoadQueue.scala 298:83:@12078.4]
  assign _T_30429 = entriesPorts_4_3 & _T_26100; // @[LoadQueue.scala 298:83:@12080.4]
  assign _T_30432 = entriesPorts_4_4 & _T_26103; // @[LoadQueue.scala 298:83:@12082.4]
  assign _T_30435 = entriesPorts_4_5 & _T_26106; // @[LoadQueue.scala 298:83:@12084.4]
  assign _T_30438 = entriesPorts_4_6 & _T_26109; // @[LoadQueue.scala 298:83:@12086.4]
  assign _T_30441 = entriesPorts_4_7 & _T_26112; // @[LoadQueue.scala 298:83:@12088.4]
  assign _T_30492 = _T_30441 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12118.4]
  assign _T_30493 = _T_30438 ? 8'h40 : _T_30492; // @[Mux.scala 31:69:@12119.4]
  assign _T_30494 = _T_30435 ? 8'h20 : _T_30493; // @[Mux.scala 31:69:@12120.4]
  assign _T_30495 = _T_30432 ? 8'h10 : _T_30494; // @[Mux.scala 31:69:@12121.4]
  assign _T_30496 = _T_30429 ? 8'h8 : _T_30495; // @[Mux.scala 31:69:@12122.4]
  assign _T_30497 = _T_30426 ? 8'h4 : _T_30496; // @[Mux.scala 31:69:@12123.4]
  assign _T_30498 = _T_30423 ? 8'h2 : _T_30497; // @[Mux.scala 31:69:@12124.4]
  assign _T_30499 = _T_30420 ? 8'h1 : _T_30498; // @[Mux.scala 31:69:@12125.4]
  assign _T_30500 = _T_30499[0]; // @[OneHot.scala 66:30:@12126.4]
  assign _T_30501 = _T_30499[1]; // @[OneHot.scala 66:30:@12127.4]
  assign _T_30502 = _T_30499[2]; // @[OneHot.scala 66:30:@12128.4]
  assign _T_30503 = _T_30499[3]; // @[OneHot.scala 66:30:@12129.4]
  assign _T_30504 = _T_30499[4]; // @[OneHot.scala 66:30:@12130.4]
  assign _T_30505 = _T_30499[5]; // @[OneHot.scala 66:30:@12131.4]
  assign _T_30506 = _T_30499[6]; // @[OneHot.scala 66:30:@12132.4]
  assign _T_30507 = _T_30499[7]; // @[OneHot.scala 66:30:@12133.4]
  assign _T_30532 = _T_30420 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12143.4]
  assign _T_30533 = _T_30441 ? 8'h40 : _T_30532; // @[Mux.scala 31:69:@12144.4]
  assign _T_30534 = _T_30438 ? 8'h20 : _T_30533; // @[Mux.scala 31:69:@12145.4]
  assign _T_30535 = _T_30435 ? 8'h10 : _T_30534; // @[Mux.scala 31:69:@12146.4]
  assign _T_30536 = _T_30432 ? 8'h8 : _T_30535; // @[Mux.scala 31:69:@12147.4]
  assign _T_30537 = _T_30429 ? 8'h4 : _T_30536; // @[Mux.scala 31:69:@12148.4]
  assign _T_30538 = _T_30426 ? 8'h2 : _T_30537; // @[Mux.scala 31:69:@12149.4]
  assign _T_30539 = _T_30423 ? 8'h1 : _T_30538; // @[Mux.scala 31:69:@12150.4]
  assign _T_30540 = _T_30539[0]; // @[OneHot.scala 66:30:@12151.4]
  assign _T_30541 = _T_30539[1]; // @[OneHot.scala 66:30:@12152.4]
  assign _T_30542 = _T_30539[2]; // @[OneHot.scala 66:30:@12153.4]
  assign _T_30543 = _T_30539[3]; // @[OneHot.scala 66:30:@12154.4]
  assign _T_30544 = _T_30539[4]; // @[OneHot.scala 66:30:@12155.4]
  assign _T_30545 = _T_30539[5]; // @[OneHot.scala 66:30:@12156.4]
  assign _T_30546 = _T_30539[6]; // @[OneHot.scala 66:30:@12157.4]
  assign _T_30547 = _T_30539[7]; // @[OneHot.scala 66:30:@12158.4]
  assign _T_30572 = _T_30423 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12168.4]
  assign _T_30573 = _T_30420 ? 8'h40 : _T_30572; // @[Mux.scala 31:69:@12169.4]
  assign _T_30574 = _T_30441 ? 8'h20 : _T_30573; // @[Mux.scala 31:69:@12170.4]
  assign _T_30575 = _T_30438 ? 8'h10 : _T_30574; // @[Mux.scala 31:69:@12171.4]
  assign _T_30576 = _T_30435 ? 8'h8 : _T_30575; // @[Mux.scala 31:69:@12172.4]
  assign _T_30577 = _T_30432 ? 8'h4 : _T_30576; // @[Mux.scala 31:69:@12173.4]
  assign _T_30578 = _T_30429 ? 8'h2 : _T_30577; // @[Mux.scala 31:69:@12174.4]
  assign _T_30579 = _T_30426 ? 8'h1 : _T_30578; // @[Mux.scala 31:69:@12175.4]
  assign _T_30580 = _T_30579[0]; // @[OneHot.scala 66:30:@12176.4]
  assign _T_30581 = _T_30579[1]; // @[OneHot.scala 66:30:@12177.4]
  assign _T_30582 = _T_30579[2]; // @[OneHot.scala 66:30:@12178.4]
  assign _T_30583 = _T_30579[3]; // @[OneHot.scala 66:30:@12179.4]
  assign _T_30584 = _T_30579[4]; // @[OneHot.scala 66:30:@12180.4]
  assign _T_30585 = _T_30579[5]; // @[OneHot.scala 66:30:@12181.4]
  assign _T_30586 = _T_30579[6]; // @[OneHot.scala 66:30:@12182.4]
  assign _T_30587 = _T_30579[7]; // @[OneHot.scala 66:30:@12183.4]
  assign _T_30612 = _T_30426 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12193.4]
  assign _T_30613 = _T_30423 ? 8'h40 : _T_30612; // @[Mux.scala 31:69:@12194.4]
  assign _T_30614 = _T_30420 ? 8'h20 : _T_30613; // @[Mux.scala 31:69:@12195.4]
  assign _T_30615 = _T_30441 ? 8'h10 : _T_30614; // @[Mux.scala 31:69:@12196.4]
  assign _T_30616 = _T_30438 ? 8'h8 : _T_30615; // @[Mux.scala 31:69:@12197.4]
  assign _T_30617 = _T_30435 ? 8'h4 : _T_30616; // @[Mux.scala 31:69:@12198.4]
  assign _T_30618 = _T_30432 ? 8'h2 : _T_30617; // @[Mux.scala 31:69:@12199.4]
  assign _T_30619 = _T_30429 ? 8'h1 : _T_30618; // @[Mux.scala 31:69:@12200.4]
  assign _T_30620 = _T_30619[0]; // @[OneHot.scala 66:30:@12201.4]
  assign _T_30621 = _T_30619[1]; // @[OneHot.scala 66:30:@12202.4]
  assign _T_30622 = _T_30619[2]; // @[OneHot.scala 66:30:@12203.4]
  assign _T_30623 = _T_30619[3]; // @[OneHot.scala 66:30:@12204.4]
  assign _T_30624 = _T_30619[4]; // @[OneHot.scala 66:30:@12205.4]
  assign _T_30625 = _T_30619[5]; // @[OneHot.scala 66:30:@12206.4]
  assign _T_30626 = _T_30619[6]; // @[OneHot.scala 66:30:@12207.4]
  assign _T_30627 = _T_30619[7]; // @[OneHot.scala 66:30:@12208.4]
  assign _T_30652 = _T_30429 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12218.4]
  assign _T_30653 = _T_30426 ? 8'h40 : _T_30652; // @[Mux.scala 31:69:@12219.4]
  assign _T_30654 = _T_30423 ? 8'h20 : _T_30653; // @[Mux.scala 31:69:@12220.4]
  assign _T_30655 = _T_30420 ? 8'h10 : _T_30654; // @[Mux.scala 31:69:@12221.4]
  assign _T_30656 = _T_30441 ? 8'h8 : _T_30655; // @[Mux.scala 31:69:@12222.4]
  assign _T_30657 = _T_30438 ? 8'h4 : _T_30656; // @[Mux.scala 31:69:@12223.4]
  assign _T_30658 = _T_30435 ? 8'h2 : _T_30657; // @[Mux.scala 31:69:@12224.4]
  assign _T_30659 = _T_30432 ? 8'h1 : _T_30658; // @[Mux.scala 31:69:@12225.4]
  assign _T_30660 = _T_30659[0]; // @[OneHot.scala 66:30:@12226.4]
  assign _T_30661 = _T_30659[1]; // @[OneHot.scala 66:30:@12227.4]
  assign _T_30662 = _T_30659[2]; // @[OneHot.scala 66:30:@12228.4]
  assign _T_30663 = _T_30659[3]; // @[OneHot.scala 66:30:@12229.4]
  assign _T_30664 = _T_30659[4]; // @[OneHot.scala 66:30:@12230.4]
  assign _T_30665 = _T_30659[5]; // @[OneHot.scala 66:30:@12231.4]
  assign _T_30666 = _T_30659[6]; // @[OneHot.scala 66:30:@12232.4]
  assign _T_30667 = _T_30659[7]; // @[OneHot.scala 66:30:@12233.4]
  assign _T_30692 = _T_30432 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12243.4]
  assign _T_30693 = _T_30429 ? 8'h40 : _T_30692; // @[Mux.scala 31:69:@12244.4]
  assign _T_30694 = _T_30426 ? 8'h20 : _T_30693; // @[Mux.scala 31:69:@12245.4]
  assign _T_30695 = _T_30423 ? 8'h10 : _T_30694; // @[Mux.scala 31:69:@12246.4]
  assign _T_30696 = _T_30420 ? 8'h8 : _T_30695; // @[Mux.scala 31:69:@12247.4]
  assign _T_30697 = _T_30441 ? 8'h4 : _T_30696; // @[Mux.scala 31:69:@12248.4]
  assign _T_30698 = _T_30438 ? 8'h2 : _T_30697; // @[Mux.scala 31:69:@12249.4]
  assign _T_30699 = _T_30435 ? 8'h1 : _T_30698; // @[Mux.scala 31:69:@12250.4]
  assign _T_30700 = _T_30699[0]; // @[OneHot.scala 66:30:@12251.4]
  assign _T_30701 = _T_30699[1]; // @[OneHot.scala 66:30:@12252.4]
  assign _T_30702 = _T_30699[2]; // @[OneHot.scala 66:30:@12253.4]
  assign _T_30703 = _T_30699[3]; // @[OneHot.scala 66:30:@12254.4]
  assign _T_30704 = _T_30699[4]; // @[OneHot.scala 66:30:@12255.4]
  assign _T_30705 = _T_30699[5]; // @[OneHot.scala 66:30:@12256.4]
  assign _T_30706 = _T_30699[6]; // @[OneHot.scala 66:30:@12257.4]
  assign _T_30707 = _T_30699[7]; // @[OneHot.scala 66:30:@12258.4]
  assign _T_30732 = _T_30435 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12268.4]
  assign _T_30733 = _T_30432 ? 8'h40 : _T_30732; // @[Mux.scala 31:69:@12269.4]
  assign _T_30734 = _T_30429 ? 8'h20 : _T_30733; // @[Mux.scala 31:69:@12270.4]
  assign _T_30735 = _T_30426 ? 8'h10 : _T_30734; // @[Mux.scala 31:69:@12271.4]
  assign _T_30736 = _T_30423 ? 8'h8 : _T_30735; // @[Mux.scala 31:69:@12272.4]
  assign _T_30737 = _T_30420 ? 8'h4 : _T_30736; // @[Mux.scala 31:69:@12273.4]
  assign _T_30738 = _T_30441 ? 8'h2 : _T_30737; // @[Mux.scala 31:69:@12274.4]
  assign _T_30739 = _T_30438 ? 8'h1 : _T_30738; // @[Mux.scala 31:69:@12275.4]
  assign _T_30740 = _T_30739[0]; // @[OneHot.scala 66:30:@12276.4]
  assign _T_30741 = _T_30739[1]; // @[OneHot.scala 66:30:@12277.4]
  assign _T_30742 = _T_30739[2]; // @[OneHot.scala 66:30:@12278.4]
  assign _T_30743 = _T_30739[3]; // @[OneHot.scala 66:30:@12279.4]
  assign _T_30744 = _T_30739[4]; // @[OneHot.scala 66:30:@12280.4]
  assign _T_30745 = _T_30739[5]; // @[OneHot.scala 66:30:@12281.4]
  assign _T_30746 = _T_30739[6]; // @[OneHot.scala 66:30:@12282.4]
  assign _T_30747 = _T_30739[7]; // @[OneHot.scala 66:30:@12283.4]
  assign _T_30772 = _T_30438 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12293.4]
  assign _T_30773 = _T_30435 ? 8'h40 : _T_30772; // @[Mux.scala 31:69:@12294.4]
  assign _T_30774 = _T_30432 ? 8'h20 : _T_30773; // @[Mux.scala 31:69:@12295.4]
  assign _T_30775 = _T_30429 ? 8'h10 : _T_30774; // @[Mux.scala 31:69:@12296.4]
  assign _T_30776 = _T_30426 ? 8'h8 : _T_30775; // @[Mux.scala 31:69:@12297.4]
  assign _T_30777 = _T_30423 ? 8'h4 : _T_30776; // @[Mux.scala 31:69:@12298.4]
  assign _T_30778 = _T_30420 ? 8'h2 : _T_30777; // @[Mux.scala 31:69:@12299.4]
  assign _T_30779 = _T_30441 ? 8'h1 : _T_30778; // @[Mux.scala 31:69:@12300.4]
  assign _T_30780 = _T_30779[0]; // @[OneHot.scala 66:30:@12301.4]
  assign _T_30781 = _T_30779[1]; // @[OneHot.scala 66:30:@12302.4]
  assign _T_30782 = _T_30779[2]; // @[OneHot.scala 66:30:@12303.4]
  assign _T_30783 = _T_30779[3]; // @[OneHot.scala 66:30:@12304.4]
  assign _T_30784 = _T_30779[4]; // @[OneHot.scala 66:30:@12305.4]
  assign _T_30785 = _T_30779[5]; // @[OneHot.scala 66:30:@12306.4]
  assign _T_30786 = _T_30779[6]; // @[OneHot.scala 66:30:@12307.4]
  assign _T_30787 = _T_30779[7]; // @[OneHot.scala 66:30:@12308.4]
  assign _T_30828 = {_T_30507,_T_30506,_T_30505,_T_30504,_T_30503,_T_30502,_T_30501,_T_30500}; // @[Mux.scala 19:72:@12324.4]
  assign _T_30830 = _T_24176 ? _T_30828 : 8'h0; // @[Mux.scala 19:72:@12325.4]
  assign _T_30837 = {_T_30546,_T_30545,_T_30544,_T_30543,_T_30542,_T_30541,_T_30540,_T_30547}; // @[Mux.scala 19:72:@12332.4]
  assign _T_30839 = _T_24177 ? _T_30837 : 8'h0; // @[Mux.scala 19:72:@12333.4]
  assign _T_30846 = {_T_30585,_T_30584,_T_30583,_T_30582,_T_30581,_T_30580,_T_30587,_T_30586}; // @[Mux.scala 19:72:@12340.4]
  assign _T_30848 = _T_24178 ? _T_30846 : 8'h0; // @[Mux.scala 19:72:@12341.4]
  assign _T_30855 = {_T_30624,_T_30623,_T_30622,_T_30621,_T_30620,_T_30627,_T_30626,_T_30625}; // @[Mux.scala 19:72:@12348.4]
  assign _T_30857 = _T_24179 ? _T_30855 : 8'h0; // @[Mux.scala 19:72:@12349.4]
  assign _T_30864 = {_T_30663,_T_30662,_T_30661,_T_30660,_T_30667,_T_30666,_T_30665,_T_30664}; // @[Mux.scala 19:72:@12356.4]
  assign _T_30866 = _T_24180 ? _T_30864 : 8'h0; // @[Mux.scala 19:72:@12357.4]
  assign _T_30873 = {_T_30702,_T_30701,_T_30700,_T_30707,_T_30706,_T_30705,_T_30704,_T_30703}; // @[Mux.scala 19:72:@12364.4]
  assign _T_30875 = _T_24181 ? _T_30873 : 8'h0; // @[Mux.scala 19:72:@12365.4]
  assign _T_30882 = {_T_30741,_T_30740,_T_30747,_T_30746,_T_30745,_T_30744,_T_30743,_T_30742}; // @[Mux.scala 19:72:@12372.4]
  assign _T_30884 = _T_24182 ? _T_30882 : 8'h0; // @[Mux.scala 19:72:@12373.4]
  assign _T_30891 = {_T_30780,_T_30787,_T_30786,_T_30785,_T_30784,_T_30783,_T_30782,_T_30781}; // @[Mux.scala 19:72:@12380.4]
  assign _T_30893 = _T_24183 ? _T_30891 : 8'h0; // @[Mux.scala 19:72:@12381.4]
  assign _T_30894 = _T_30830 | _T_30839; // @[Mux.scala 19:72:@12382.4]
  assign _T_30895 = _T_30894 | _T_30848; // @[Mux.scala 19:72:@12383.4]
  assign _T_30896 = _T_30895 | _T_30857; // @[Mux.scala 19:72:@12384.4]
  assign _T_30897 = _T_30896 | _T_30866; // @[Mux.scala 19:72:@12385.4]
  assign _T_30898 = _T_30897 | _T_30875; // @[Mux.scala 19:72:@12386.4]
  assign _T_30899 = _T_30898 | _T_30884; // @[Mux.scala 19:72:@12387.4]
  assign _T_30900 = _T_30899 | _T_30893; // @[Mux.scala 19:72:@12388.4]
  assign inputPriorityPorts_4_0 = _T_30900[0]; // @[Mux.scala 19:72:@12392.4]
  assign inputPriorityPorts_4_1 = _T_30900[1]; // @[Mux.scala 19:72:@12394.4]
  assign inputPriorityPorts_4_2 = _T_30900[2]; // @[Mux.scala 19:72:@12396.4]
  assign inputPriorityPorts_4_3 = _T_30900[3]; // @[Mux.scala 19:72:@12398.4]
  assign inputPriorityPorts_4_4 = _T_30900[4]; // @[Mux.scala 19:72:@12400.4]
  assign inputPriorityPorts_4_5 = _T_30900[5]; // @[Mux.scala 19:72:@12402.4]
  assign inputPriorityPorts_4_6 = _T_30900[6]; // @[Mux.scala 19:72:@12404.4]
  assign inputPriorityPorts_4_7 = _T_30900[7]; // @[Mux.scala 19:72:@12406.4]
  assign _T_31014 = entriesPorts_4_7 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12436.4]
  assign _T_31015 = entriesPorts_4_6 ? 8'h40 : _T_31014; // @[Mux.scala 31:69:@12437.4]
  assign _T_31016 = entriesPorts_4_5 ? 8'h20 : _T_31015; // @[Mux.scala 31:69:@12438.4]
  assign _T_31017 = entriesPorts_4_4 ? 8'h10 : _T_31016; // @[Mux.scala 31:69:@12439.4]
  assign _T_31018 = entriesPorts_4_3 ? 8'h8 : _T_31017; // @[Mux.scala 31:69:@12440.4]
  assign _T_31019 = entriesPorts_4_2 ? 8'h4 : _T_31018; // @[Mux.scala 31:69:@12441.4]
  assign _T_31020 = entriesPorts_4_1 ? 8'h2 : _T_31019; // @[Mux.scala 31:69:@12442.4]
  assign _T_31021 = entriesPorts_4_0 ? 8'h1 : _T_31020; // @[Mux.scala 31:69:@12443.4]
  assign _T_31022 = _T_31021[0]; // @[OneHot.scala 66:30:@12444.4]
  assign _T_31023 = _T_31021[1]; // @[OneHot.scala 66:30:@12445.4]
  assign _T_31024 = _T_31021[2]; // @[OneHot.scala 66:30:@12446.4]
  assign _T_31025 = _T_31021[3]; // @[OneHot.scala 66:30:@12447.4]
  assign _T_31026 = _T_31021[4]; // @[OneHot.scala 66:30:@12448.4]
  assign _T_31027 = _T_31021[5]; // @[OneHot.scala 66:30:@12449.4]
  assign _T_31028 = _T_31021[6]; // @[OneHot.scala 66:30:@12450.4]
  assign _T_31029 = _T_31021[7]; // @[OneHot.scala 66:30:@12451.4]
  assign _T_31054 = entriesPorts_4_0 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12461.4]
  assign _T_31055 = entriesPorts_4_7 ? 8'h40 : _T_31054; // @[Mux.scala 31:69:@12462.4]
  assign _T_31056 = entriesPorts_4_6 ? 8'h20 : _T_31055; // @[Mux.scala 31:69:@12463.4]
  assign _T_31057 = entriesPorts_4_5 ? 8'h10 : _T_31056; // @[Mux.scala 31:69:@12464.4]
  assign _T_31058 = entriesPorts_4_4 ? 8'h8 : _T_31057; // @[Mux.scala 31:69:@12465.4]
  assign _T_31059 = entriesPorts_4_3 ? 8'h4 : _T_31058; // @[Mux.scala 31:69:@12466.4]
  assign _T_31060 = entriesPorts_4_2 ? 8'h2 : _T_31059; // @[Mux.scala 31:69:@12467.4]
  assign _T_31061 = entriesPorts_4_1 ? 8'h1 : _T_31060; // @[Mux.scala 31:69:@12468.4]
  assign _T_31062 = _T_31061[0]; // @[OneHot.scala 66:30:@12469.4]
  assign _T_31063 = _T_31061[1]; // @[OneHot.scala 66:30:@12470.4]
  assign _T_31064 = _T_31061[2]; // @[OneHot.scala 66:30:@12471.4]
  assign _T_31065 = _T_31061[3]; // @[OneHot.scala 66:30:@12472.4]
  assign _T_31066 = _T_31061[4]; // @[OneHot.scala 66:30:@12473.4]
  assign _T_31067 = _T_31061[5]; // @[OneHot.scala 66:30:@12474.4]
  assign _T_31068 = _T_31061[6]; // @[OneHot.scala 66:30:@12475.4]
  assign _T_31069 = _T_31061[7]; // @[OneHot.scala 66:30:@12476.4]
  assign _T_31094 = entriesPorts_4_1 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12486.4]
  assign _T_31095 = entriesPorts_4_0 ? 8'h40 : _T_31094; // @[Mux.scala 31:69:@12487.4]
  assign _T_31096 = entriesPorts_4_7 ? 8'h20 : _T_31095; // @[Mux.scala 31:69:@12488.4]
  assign _T_31097 = entriesPorts_4_6 ? 8'h10 : _T_31096; // @[Mux.scala 31:69:@12489.4]
  assign _T_31098 = entriesPorts_4_5 ? 8'h8 : _T_31097; // @[Mux.scala 31:69:@12490.4]
  assign _T_31099 = entriesPorts_4_4 ? 8'h4 : _T_31098; // @[Mux.scala 31:69:@12491.4]
  assign _T_31100 = entriesPorts_4_3 ? 8'h2 : _T_31099; // @[Mux.scala 31:69:@12492.4]
  assign _T_31101 = entriesPorts_4_2 ? 8'h1 : _T_31100; // @[Mux.scala 31:69:@12493.4]
  assign _T_31102 = _T_31101[0]; // @[OneHot.scala 66:30:@12494.4]
  assign _T_31103 = _T_31101[1]; // @[OneHot.scala 66:30:@12495.4]
  assign _T_31104 = _T_31101[2]; // @[OneHot.scala 66:30:@12496.4]
  assign _T_31105 = _T_31101[3]; // @[OneHot.scala 66:30:@12497.4]
  assign _T_31106 = _T_31101[4]; // @[OneHot.scala 66:30:@12498.4]
  assign _T_31107 = _T_31101[5]; // @[OneHot.scala 66:30:@12499.4]
  assign _T_31108 = _T_31101[6]; // @[OneHot.scala 66:30:@12500.4]
  assign _T_31109 = _T_31101[7]; // @[OneHot.scala 66:30:@12501.4]
  assign _T_31134 = entriesPorts_4_2 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12511.4]
  assign _T_31135 = entriesPorts_4_1 ? 8'h40 : _T_31134; // @[Mux.scala 31:69:@12512.4]
  assign _T_31136 = entriesPorts_4_0 ? 8'h20 : _T_31135; // @[Mux.scala 31:69:@12513.4]
  assign _T_31137 = entriesPorts_4_7 ? 8'h10 : _T_31136; // @[Mux.scala 31:69:@12514.4]
  assign _T_31138 = entriesPorts_4_6 ? 8'h8 : _T_31137; // @[Mux.scala 31:69:@12515.4]
  assign _T_31139 = entriesPorts_4_5 ? 8'h4 : _T_31138; // @[Mux.scala 31:69:@12516.4]
  assign _T_31140 = entriesPorts_4_4 ? 8'h2 : _T_31139; // @[Mux.scala 31:69:@12517.4]
  assign _T_31141 = entriesPorts_4_3 ? 8'h1 : _T_31140; // @[Mux.scala 31:69:@12518.4]
  assign _T_31142 = _T_31141[0]; // @[OneHot.scala 66:30:@12519.4]
  assign _T_31143 = _T_31141[1]; // @[OneHot.scala 66:30:@12520.4]
  assign _T_31144 = _T_31141[2]; // @[OneHot.scala 66:30:@12521.4]
  assign _T_31145 = _T_31141[3]; // @[OneHot.scala 66:30:@12522.4]
  assign _T_31146 = _T_31141[4]; // @[OneHot.scala 66:30:@12523.4]
  assign _T_31147 = _T_31141[5]; // @[OneHot.scala 66:30:@12524.4]
  assign _T_31148 = _T_31141[6]; // @[OneHot.scala 66:30:@12525.4]
  assign _T_31149 = _T_31141[7]; // @[OneHot.scala 66:30:@12526.4]
  assign _T_31174 = entriesPorts_4_3 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12536.4]
  assign _T_31175 = entriesPorts_4_2 ? 8'h40 : _T_31174; // @[Mux.scala 31:69:@12537.4]
  assign _T_31176 = entriesPorts_4_1 ? 8'h20 : _T_31175; // @[Mux.scala 31:69:@12538.4]
  assign _T_31177 = entriesPorts_4_0 ? 8'h10 : _T_31176; // @[Mux.scala 31:69:@12539.4]
  assign _T_31178 = entriesPorts_4_7 ? 8'h8 : _T_31177; // @[Mux.scala 31:69:@12540.4]
  assign _T_31179 = entriesPorts_4_6 ? 8'h4 : _T_31178; // @[Mux.scala 31:69:@12541.4]
  assign _T_31180 = entriesPorts_4_5 ? 8'h2 : _T_31179; // @[Mux.scala 31:69:@12542.4]
  assign _T_31181 = entriesPorts_4_4 ? 8'h1 : _T_31180; // @[Mux.scala 31:69:@12543.4]
  assign _T_31182 = _T_31181[0]; // @[OneHot.scala 66:30:@12544.4]
  assign _T_31183 = _T_31181[1]; // @[OneHot.scala 66:30:@12545.4]
  assign _T_31184 = _T_31181[2]; // @[OneHot.scala 66:30:@12546.4]
  assign _T_31185 = _T_31181[3]; // @[OneHot.scala 66:30:@12547.4]
  assign _T_31186 = _T_31181[4]; // @[OneHot.scala 66:30:@12548.4]
  assign _T_31187 = _T_31181[5]; // @[OneHot.scala 66:30:@12549.4]
  assign _T_31188 = _T_31181[6]; // @[OneHot.scala 66:30:@12550.4]
  assign _T_31189 = _T_31181[7]; // @[OneHot.scala 66:30:@12551.4]
  assign _T_31214 = entriesPorts_4_4 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12561.4]
  assign _T_31215 = entriesPorts_4_3 ? 8'h40 : _T_31214; // @[Mux.scala 31:69:@12562.4]
  assign _T_31216 = entriesPorts_4_2 ? 8'h20 : _T_31215; // @[Mux.scala 31:69:@12563.4]
  assign _T_31217 = entriesPorts_4_1 ? 8'h10 : _T_31216; // @[Mux.scala 31:69:@12564.4]
  assign _T_31218 = entriesPorts_4_0 ? 8'h8 : _T_31217; // @[Mux.scala 31:69:@12565.4]
  assign _T_31219 = entriesPorts_4_7 ? 8'h4 : _T_31218; // @[Mux.scala 31:69:@12566.4]
  assign _T_31220 = entriesPorts_4_6 ? 8'h2 : _T_31219; // @[Mux.scala 31:69:@12567.4]
  assign _T_31221 = entriesPorts_4_5 ? 8'h1 : _T_31220; // @[Mux.scala 31:69:@12568.4]
  assign _T_31222 = _T_31221[0]; // @[OneHot.scala 66:30:@12569.4]
  assign _T_31223 = _T_31221[1]; // @[OneHot.scala 66:30:@12570.4]
  assign _T_31224 = _T_31221[2]; // @[OneHot.scala 66:30:@12571.4]
  assign _T_31225 = _T_31221[3]; // @[OneHot.scala 66:30:@12572.4]
  assign _T_31226 = _T_31221[4]; // @[OneHot.scala 66:30:@12573.4]
  assign _T_31227 = _T_31221[5]; // @[OneHot.scala 66:30:@12574.4]
  assign _T_31228 = _T_31221[6]; // @[OneHot.scala 66:30:@12575.4]
  assign _T_31229 = _T_31221[7]; // @[OneHot.scala 66:30:@12576.4]
  assign _T_31254 = entriesPorts_4_5 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12586.4]
  assign _T_31255 = entriesPorts_4_4 ? 8'h40 : _T_31254; // @[Mux.scala 31:69:@12587.4]
  assign _T_31256 = entriesPorts_4_3 ? 8'h20 : _T_31255; // @[Mux.scala 31:69:@12588.4]
  assign _T_31257 = entriesPorts_4_2 ? 8'h10 : _T_31256; // @[Mux.scala 31:69:@12589.4]
  assign _T_31258 = entriesPorts_4_1 ? 8'h8 : _T_31257; // @[Mux.scala 31:69:@12590.4]
  assign _T_31259 = entriesPorts_4_0 ? 8'h4 : _T_31258; // @[Mux.scala 31:69:@12591.4]
  assign _T_31260 = entriesPorts_4_7 ? 8'h2 : _T_31259; // @[Mux.scala 31:69:@12592.4]
  assign _T_31261 = entriesPorts_4_6 ? 8'h1 : _T_31260; // @[Mux.scala 31:69:@12593.4]
  assign _T_31262 = _T_31261[0]; // @[OneHot.scala 66:30:@12594.4]
  assign _T_31263 = _T_31261[1]; // @[OneHot.scala 66:30:@12595.4]
  assign _T_31264 = _T_31261[2]; // @[OneHot.scala 66:30:@12596.4]
  assign _T_31265 = _T_31261[3]; // @[OneHot.scala 66:30:@12597.4]
  assign _T_31266 = _T_31261[4]; // @[OneHot.scala 66:30:@12598.4]
  assign _T_31267 = _T_31261[5]; // @[OneHot.scala 66:30:@12599.4]
  assign _T_31268 = _T_31261[6]; // @[OneHot.scala 66:30:@12600.4]
  assign _T_31269 = _T_31261[7]; // @[OneHot.scala 66:30:@12601.4]
  assign _T_31294 = entriesPorts_4_6 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@12611.4]
  assign _T_31295 = entriesPorts_4_5 ? 8'h40 : _T_31294; // @[Mux.scala 31:69:@12612.4]
  assign _T_31296 = entriesPorts_4_4 ? 8'h20 : _T_31295; // @[Mux.scala 31:69:@12613.4]
  assign _T_31297 = entriesPorts_4_3 ? 8'h10 : _T_31296; // @[Mux.scala 31:69:@12614.4]
  assign _T_31298 = entriesPorts_4_2 ? 8'h8 : _T_31297; // @[Mux.scala 31:69:@12615.4]
  assign _T_31299 = entriesPorts_4_1 ? 8'h4 : _T_31298; // @[Mux.scala 31:69:@12616.4]
  assign _T_31300 = entriesPorts_4_0 ? 8'h2 : _T_31299; // @[Mux.scala 31:69:@12617.4]
  assign _T_31301 = entriesPorts_4_7 ? 8'h1 : _T_31300; // @[Mux.scala 31:69:@12618.4]
  assign _T_31302 = _T_31301[0]; // @[OneHot.scala 66:30:@12619.4]
  assign _T_31303 = _T_31301[1]; // @[OneHot.scala 66:30:@12620.4]
  assign _T_31304 = _T_31301[2]; // @[OneHot.scala 66:30:@12621.4]
  assign _T_31305 = _T_31301[3]; // @[OneHot.scala 66:30:@12622.4]
  assign _T_31306 = _T_31301[4]; // @[OneHot.scala 66:30:@12623.4]
  assign _T_31307 = _T_31301[5]; // @[OneHot.scala 66:30:@12624.4]
  assign _T_31308 = _T_31301[6]; // @[OneHot.scala 66:30:@12625.4]
  assign _T_31309 = _T_31301[7]; // @[OneHot.scala 66:30:@12626.4]
  assign _T_31350 = {_T_31029,_T_31028,_T_31027,_T_31026,_T_31025,_T_31024,_T_31023,_T_31022}; // @[Mux.scala 19:72:@12642.4]
  assign _T_31352 = _T_24176 ? _T_31350 : 8'h0; // @[Mux.scala 19:72:@12643.4]
  assign _T_31359 = {_T_31068,_T_31067,_T_31066,_T_31065,_T_31064,_T_31063,_T_31062,_T_31069}; // @[Mux.scala 19:72:@12650.4]
  assign _T_31361 = _T_24177 ? _T_31359 : 8'h0; // @[Mux.scala 19:72:@12651.4]
  assign _T_31368 = {_T_31107,_T_31106,_T_31105,_T_31104,_T_31103,_T_31102,_T_31109,_T_31108}; // @[Mux.scala 19:72:@12658.4]
  assign _T_31370 = _T_24178 ? _T_31368 : 8'h0; // @[Mux.scala 19:72:@12659.4]
  assign _T_31377 = {_T_31146,_T_31145,_T_31144,_T_31143,_T_31142,_T_31149,_T_31148,_T_31147}; // @[Mux.scala 19:72:@12666.4]
  assign _T_31379 = _T_24179 ? _T_31377 : 8'h0; // @[Mux.scala 19:72:@12667.4]
  assign _T_31386 = {_T_31185,_T_31184,_T_31183,_T_31182,_T_31189,_T_31188,_T_31187,_T_31186}; // @[Mux.scala 19:72:@12674.4]
  assign _T_31388 = _T_24180 ? _T_31386 : 8'h0; // @[Mux.scala 19:72:@12675.4]
  assign _T_31395 = {_T_31224,_T_31223,_T_31222,_T_31229,_T_31228,_T_31227,_T_31226,_T_31225}; // @[Mux.scala 19:72:@12682.4]
  assign _T_31397 = _T_24181 ? _T_31395 : 8'h0; // @[Mux.scala 19:72:@12683.4]
  assign _T_31404 = {_T_31263,_T_31262,_T_31269,_T_31268,_T_31267,_T_31266,_T_31265,_T_31264}; // @[Mux.scala 19:72:@12690.4]
  assign _T_31406 = _T_24182 ? _T_31404 : 8'h0; // @[Mux.scala 19:72:@12691.4]
  assign _T_31413 = {_T_31302,_T_31309,_T_31308,_T_31307,_T_31306,_T_31305,_T_31304,_T_31303}; // @[Mux.scala 19:72:@12698.4]
  assign _T_31415 = _T_24183 ? _T_31413 : 8'h0; // @[Mux.scala 19:72:@12699.4]
  assign _T_31416 = _T_31352 | _T_31361; // @[Mux.scala 19:72:@12700.4]
  assign _T_31417 = _T_31416 | _T_31370; // @[Mux.scala 19:72:@12701.4]
  assign _T_31418 = _T_31417 | _T_31379; // @[Mux.scala 19:72:@12702.4]
  assign _T_31419 = _T_31418 | _T_31388; // @[Mux.scala 19:72:@12703.4]
  assign _T_31420 = _T_31419 | _T_31397; // @[Mux.scala 19:72:@12704.4]
  assign _T_31421 = _T_31420 | _T_31406; // @[Mux.scala 19:72:@12705.4]
  assign _T_31422 = _T_31421 | _T_31415; // @[Mux.scala 19:72:@12706.4]
  assign outputPriorityPorts_4_0 = _T_31422[0]; // @[Mux.scala 19:72:@12710.4]
  assign outputPriorityPorts_4_1 = _T_31422[1]; // @[Mux.scala 19:72:@12712.4]
  assign outputPriorityPorts_4_2 = _T_31422[2]; // @[Mux.scala 19:72:@12714.4]
  assign outputPriorityPorts_4_3 = _T_31422[3]; // @[Mux.scala 19:72:@12716.4]
  assign outputPriorityPorts_4_4 = _T_31422[4]; // @[Mux.scala 19:72:@12718.4]
  assign outputPriorityPorts_4_5 = _T_31422[5]; // @[Mux.scala 19:72:@12720.4]
  assign outputPriorityPorts_4_6 = _T_31422[6]; // @[Mux.scala 19:72:@12722.4]
  assign outputPriorityPorts_4_7 = _T_31422[7]; // @[Mux.scala 19:72:@12724.4]
  assign _T_31501 = inputPriorityPorts_0_0 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@12738.6]
  assign _T_31502 = inputPriorityPorts_1_0 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@12739.6]
  assign _T_31503 = inputPriorityPorts_2_0 & io_loadAddrEnable_2; // @[LoadQueue.scala 313:47:@12740.6]
  assign _T_31504 = inputPriorityPorts_3_0 & io_loadAddrEnable_3; // @[LoadQueue.scala 313:47:@12741.6]
  assign _T_31505 = inputPriorityPorts_4_0 & io_loadAddrEnable_4; // @[LoadQueue.scala 313:47:@12742.6]
  assign _T_31519 = _T_31501 | _T_31502; // @[LoadQueue.scala 314:26:@12750.6]
  assign _T_31520 = _T_31519 | _T_31503; // @[LoadQueue.scala 314:26:@12751.6]
  assign _T_31521 = _T_31520 | _T_31504; // @[LoadQueue.scala 314:26:@12752.6]
  assign _T_31522 = _T_31521 | _T_31505; // @[LoadQueue.scala 314:26:@12753.6]
  assign _T_31526 = {_T_31505,_T_31504,_T_31503,_T_31502,_T_31501}; // @[OneHot.scala 18:45:@12758.8]
  assign _T_31527 = _T_31526[4]; // @[OneHot.scala 26:18:@12759.8]
  assign _T_31528 = _T_31526[3:0]; // @[OneHot.scala 27:18:@12760.8]
  assign _GEN_814 = {{3'd0}, _T_31527}; // @[OneHot.scala 28:28:@12762.8]
  assign _T_31531 = _GEN_814 | _T_31528; // @[OneHot.scala 28:28:@12762.8]
  assign _T_31532 = _T_31531[3:2]; // @[OneHot.scala 26:18:@12763.8]
  assign _T_31533 = _T_31531[1:0]; // @[OneHot.scala 27:18:@12764.8]
  assign _T_31535 = _T_31532 != 2'h0; // @[OneHot.scala 28:14:@12765.8]
  assign _T_31536 = _T_31532 | _T_31533; // @[OneHot.scala 28:28:@12766.8]
  assign _T_31537 = _T_31536[1]; // @[CircuitMath.scala 30:8:@12767.8]
  assign _T_31539 = {_T_31527,_T_31535,_T_31537}; // @[Cat.scala 30:58:@12769.8]
  assign _GEN_611 = 3'h1 == _T_31539 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@12770.8]
  assign _GEN_612 = 3'h2 == _T_31539 ? io_addrFromLoadPorts_2 : _GEN_611; // @[LoadQueue.scala 315:29:@12770.8]
  assign _GEN_613 = 3'h3 == _T_31539 ? io_addrFromLoadPorts_3 : _GEN_612; // @[LoadQueue.scala 315:29:@12770.8]
  assign _GEN_614 = 3'h4 == _T_31539 ? io_addrFromLoadPorts_4 : _GEN_613; // @[LoadQueue.scala 315:29:@12770.8]
  assign _GEN_615 = _T_31522 ? _GEN_614 : addrQ_0; // @[LoadQueue.scala 314:36:@12754.6]
  assign _GEN_616 = _T_31522 ? 1'h1 : addrKnown_0; // @[LoadQueue.scala 314:36:@12754.6]
  assign _GEN_617 = initBits_0 ? 1'h0 : _GEN_616; // @[LoadQueue.scala 308:34:@12734.4]
  assign _GEN_618 = initBits_0 ? addrQ_0 : _GEN_615; // @[LoadQueue.scala 308:34:@12734.4]
  assign _T_31543 = inputPriorityPorts_0_1 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@12778.6]
  assign _T_31544 = inputPriorityPorts_1_1 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@12779.6]
  assign _T_31545 = inputPriorityPorts_2_1 & io_loadAddrEnable_2; // @[LoadQueue.scala 313:47:@12780.6]
  assign _T_31546 = inputPriorityPorts_3_1 & io_loadAddrEnable_3; // @[LoadQueue.scala 313:47:@12781.6]
  assign _T_31547 = inputPriorityPorts_4_1 & io_loadAddrEnable_4; // @[LoadQueue.scala 313:47:@12782.6]
  assign _T_31561 = _T_31543 | _T_31544; // @[LoadQueue.scala 314:26:@12790.6]
  assign _T_31562 = _T_31561 | _T_31545; // @[LoadQueue.scala 314:26:@12791.6]
  assign _T_31563 = _T_31562 | _T_31546; // @[LoadQueue.scala 314:26:@12792.6]
  assign _T_31564 = _T_31563 | _T_31547; // @[LoadQueue.scala 314:26:@12793.6]
  assign _T_31568 = {_T_31547,_T_31546,_T_31545,_T_31544,_T_31543}; // @[OneHot.scala 18:45:@12798.8]
  assign _T_31569 = _T_31568[4]; // @[OneHot.scala 26:18:@12799.8]
  assign _T_31570 = _T_31568[3:0]; // @[OneHot.scala 27:18:@12800.8]
  assign _GEN_815 = {{3'd0}, _T_31569}; // @[OneHot.scala 28:28:@12802.8]
  assign _T_31573 = _GEN_815 | _T_31570; // @[OneHot.scala 28:28:@12802.8]
  assign _T_31574 = _T_31573[3:2]; // @[OneHot.scala 26:18:@12803.8]
  assign _T_31575 = _T_31573[1:0]; // @[OneHot.scala 27:18:@12804.8]
  assign _T_31577 = _T_31574 != 2'h0; // @[OneHot.scala 28:14:@12805.8]
  assign _T_31578 = _T_31574 | _T_31575; // @[OneHot.scala 28:28:@12806.8]
  assign _T_31579 = _T_31578[1]; // @[CircuitMath.scala 30:8:@12807.8]
  assign _T_31581 = {_T_31569,_T_31577,_T_31579}; // @[Cat.scala 30:58:@12809.8]
  assign _GEN_620 = 3'h1 == _T_31581 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@12810.8]
  assign _GEN_621 = 3'h2 == _T_31581 ? io_addrFromLoadPorts_2 : _GEN_620; // @[LoadQueue.scala 315:29:@12810.8]
  assign _GEN_622 = 3'h3 == _T_31581 ? io_addrFromLoadPorts_3 : _GEN_621; // @[LoadQueue.scala 315:29:@12810.8]
  assign _GEN_623 = 3'h4 == _T_31581 ? io_addrFromLoadPorts_4 : _GEN_622; // @[LoadQueue.scala 315:29:@12810.8]
  assign _GEN_624 = _T_31564 ? _GEN_623 : addrQ_1; // @[LoadQueue.scala 314:36:@12794.6]
  assign _GEN_625 = _T_31564 ? 1'h1 : addrKnown_1; // @[LoadQueue.scala 314:36:@12794.6]
  assign _GEN_626 = initBits_1 ? 1'h0 : _GEN_625; // @[LoadQueue.scala 308:34:@12774.4]
  assign _GEN_627 = initBits_1 ? addrQ_1 : _GEN_624; // @[LoadQueue.scala 308:34:@12774.4]
  assign _T_31585 = inputPriorityPorts_0_2 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@12818.6]
  assign _T_31586 = inputPriorityPorts_1_2 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@12819.6]
  assign _T_31587 = inputPriorityPorts_2_2 & io_loadAddrEnable_2; // @[LoadQueue.scala 313:47:@12820.6]
  assign _T_31588 = inputPriorityPorts_3_2 & io_loadAddrEnable_3; // @[LoadQueue.scala 313:47:@12821.6]
  assign _T_31589 = inputPriorityPorts_4_2 & io_loadAddrEnable_4; // @[LoadQueue.scala 313:47:@12822.6]
  assign _T_31603 = _T_31585 | _T_31586; // @[LoadQueue.scala 314:26:@12830.6]
  assign _T_31604 = _T_31603 | _T_31587; // @[LoadQueue.scala 314:26:@12831.6]
  assign _T_31605 = _T_31604 | _T_31588; // @[LoadQueue.scala 314:26:@12832.6]
  assign _T_31606 = _T_31605 | _T_31589; // @[LoadQueue.scala 314:26:@12833.6]
  assign _T_31610 = {_T_31589,_T_31588,_T_31587,_T_31586,_T_31585}; // @[OneHot.scala 18:45:@12838.8]
  assign _T_31611 = _T_31610[4]; // @[OneHot.scala 26:18:@12839.8]
  assign _T_31612 = _T_31610[3:0]; // @[OneHot.scala 27:18:@12840.8]
  assign _GEN_816 = {{3'd0}, _T_31611}; // @[OneHot.scala 28:28:@12842.8]
  assign _T_31615 = _GEN_816 | _T_31612; // @[OneHot.scala 28:28:@12842.8]
  assign _T_31616 = _T_31615[3:2]; // @[OneHot.scala 26:18:@12843.8]
  assign _T_31617 = _T_31615[1:0]; // @[OneHot.scala 27:18:@12844.8]
  assign _T_31619 = _T_31616 != 2'h0; // @[OneHot.scala 28:14:@12845.8]
  assign _T_31620 = _T_31616 | _T_31617; // @[OneHot.scala 28:28:@12846.8]
  assign _T_31621 = _T_31620[1]; // @[CircuitMath.scala 30:8:@12847.8]
  assign _T_31623 = {_T_31611,_T_31619,_T_31621}; // @[Cat.scala 30:58:@12849.8]
  assign _GEN_629 = 3'h1 == _T_31623 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@12850.8]
  assign _GEN_630 = 3'h2 == _T_31623 ? io_addrFromLoadPorts_2 : _GEN_629; // @[LoadQueue.scala 315:29:@12850.8]
  assign _GEN_631 = 3'h3 == _T_31623 ? io_addrFromLoadPorts_3 : _GEN_630; // @[LoadQueue.scala 315:29:@12850.8]
  assign _GEN_632 = 3'h4 == _T_31623 ? io_addrFromLoadPorts_4 : _GEN_631; // @[LoadQueue.scala 315:29:@12850.8]
  assign _GEN_633 = _T_31606 ? _GEN_632 : addrQ_2; // @[LoadQueue.scala 314:36:@12834.6]
  assign _GEN_634 = _T_31606 ? 1'h1 : addrKnown_2; // @[LoadQueue.scala 314:36:@12834.6]
  assign _GEN_635 = initBits_2 ? 1'h0 : _GEN_634; // @[LoadQueue.scala 308:34:@12814.4]
  assign _GEN_636 = initBits_2 ? addrQ_2 : _GEN_633; // @[LoadQueue.scala 308:34:@12814.4]
  assign _T_31627 = inputPriorityPorts_0_3 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@12858.6]
  assign _T_31628 = inputPriorityPorts_1_3 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@12859.6]
  assign _T_31629 = inputPriorityPorts_2_3 & io_loadAddrEnable_2; // @[LoadQueue.scala 313:47:@12860.6]
  assign _T_31630 = inputPriorityPorts_3_3 & io_loadAddrEnable_3; // @[LoadQueue.scala 313:47:@12861.6]
  assign _T_31631 = inputPriorityPorts_4_3 & io_loadAddrEnable_4; // @[LoadQueue.scala 313:47:@12862.6]
  assign _T_31645 = _T_31627 | _T_31628; // @[LoadQueue.scala 314:26:@12870.6]
  assign _T_31646 = _T_31645 | _T_31629; // @[LoadQueue.scala 314:26:@12871.6]
  assign _T_31647 = _T_31646 | _T_31630; // @[LoadQueue.scala 314:26:@12872.6]
  assign _T_31648 = _T_31647 | _T_31631; // @[LoadQueue.scala 314:26:@12873.6]
  assign _T_31652 = {_T_31631,_T_31630,_T_31629,_T_31628,_T_31627}; // @[OneHot.scala 18:45:@12878.8]
  assign _T_31653 = _T_31652[4]; // @[OneHot.scala 26:18:@12879.8]
  assign _T_31654 = _T_31652[3:0]; // @[OneHot.scala 27:18:@12880.8]
  assign _GEN_817 = {{3'd0}, _T_31653}; // @[OneHot.scala 28:28:@12882.8]
  assign _T_31657 = _GEN_817 | _T_31654; // @[OneHot.scala 28:28:@12882.8]
  assign _T_31658 = _T_31657[3:2]; // @[OneHot.scala 26:18:@12883.8]
  assign _T_31659 = _T_31657[1:0]; // @[OneHot.scala 27:18:@12884.8]
  assign _T_31661 = _T_31658 != 2'h0; // @[OneHot.scala 28:14:@12885.8]
  assign _T_31662 = _T_31658 | _T_31659; // @[OneHot.scala 28:28:@12886.8]
  assign _T_31663 = _T_31662[1]; // @[CircuitMath.scala 30:8:@12887.8]
  assign _T_31665 = {_T_31653,_T_31661,_T_31663}; // @[Cat.scala 30:58:@12889.8]
  assign _GEN_638 = 3'h1 == _T_31665 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@12890.8]
  assign _GEN_639 = 3'h2 == _T_31665 ? io_addrFromLoadPorts_2 : _GEN_638; // @[LoadQueue.scala 315:29:@12890.8]
  assign _GEN_640 = 3'h3 == _T_31665 ? io_addrFromLoadPorts_3 : _GEN_639; // @[LoadQueue.scala 315:29:@12890.8]
  assign _GEN_641 = 3'h4 == _T_31665 ? io_addrFromLoadPorts_4 : _GEN_640; // @[LoadQueue.scala 315:29:@12890.8]
  assign _GEN_642 = _T_31648 ? _GEN_641 : addrQ_3; // @[LoadQueue.scala 314:36:@12874.6]
  assign _GEN_643 = _T_31648 ? 1'h1 : addrKnown_3; // @[LoadQueue.scala 314:36:@12874.6]
  assign _GEN_644 = initBits_3 ? 1'h0 : _GEN_643; // @[LoadQueue.scala 308:34:@12854.4]
  assign _GEN_645 = initBits_3 ? addrQ_3 : _GEN_642; // @[LoadQueue.scala 308:34:@12854.4]
  assign _T_31669 = inputPriorityPorts_0_4 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@12898.6]
  assign _T_31670 = inputPriorityPorts_1_4 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@12899.6]
  assign _T_31671 = inputPriorityPorts_2_4 & io_loadAddrEnable_2; // @[LoadQueue.scala 313:47:@12900.6]
  assign _T_31672 = inputPriorityPorts_3_4 & io_loadAddrEnable_3; // @[LoadQueue.scala 313:47:@12901.6]
  assign _T_31673 = inputPriorityPorts_4_4 & io_loadAddrEnable_4; // @[LoadQueue.scala 313:47:@12902.6]
  assign _T_31687 = _T_31669 | _T_31670; // @[LoadQueue.scala 314:26:@12910.6]
  assign _T_31688 = _T_31687 | _T_31671; // @[LoadQueue.scala 314:26:@12911.6]
  assign _T_31689 = _T_31688 | _T_31672; // @[LoadQueue.scala 314:26:@12912.6]
  assign _T_31690 = _T_31689 | _T_31673; // @[LoadQueue.scala 314:26:@12913.6]
  assign _T_31694 = {_T_31673,_T_31672,_T_31671,_T_31670,_T_31669}; // @[OneHot.scala 18:45:@12918.8]
  assign _T_31695 = _T_31694[4]; // @[OneHot.scala 26:18:@12919.8]
  assign _T_31696 = _T_31694[3:0]; // @[OneHot.scala 27:18:@12920.8]
  assign _GEN_818 = {{3'd0}, _T_31695}; // @[OneHot.scala 28:28:@12922.8]
  assign _T_31699 = _GEN_818 | _T_31696; // @[OneHot.scala 28:28:@12922.8]
  assign _T_31700 = _T_31699[3:2]; // @[OneHot.scala 26:18:@12923.8]
  assign _T_31701 = _T_31699[1:0]; // @[OneHot.scala 27:18:@12924.8]
  assign _T_31703 = _T_31700 != 2'h0; // @[OneHot.scala 28:14:@12925.8]
  assign _T_31704 = _T_31700 | _T_31701; // @[OneHot.scala 28:28:@12926.8]
  assign _T_31705 = _T_31704[1]; // @[CircuitMath.scala 30:8:@12927.8]
  assign _T_31707 = {_T_31695,_T_31703,_T_31705}; // @[Cat.scala 30:58:@12929.8]
  assign _GEN_647 = 3'h1 == _T_31707 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@12930.8]
  assign _GEN_648 = 3'h2 == _T_31707 ? io_addrFromLoadPorts_2 : _GEN_647; // @[LoadQueue.scala 315:29:@12930.8]
  assign _GEN_649 = 3'h3 == _T_31707 ? io_addrFromLoadPorts_3 : _GEN_648; // @[LoadQueue.scala 315:29:@12930.8]
  assign _GEN_650 = 3'h4 == _T_31707 ? io_addrFromLoadPorts_4 : _GEN_649; // @[LoadQueue.scala 315:29:@12930.8]
  assign _GEN_651 = _T_31690 ? _GEN_650 : addrQ_4; // @[LoadQueue.scala 314:36:@12914.6]
  assign _GEN_652 = _T_31690 ? 1'h1 : addrKnown_4; // @[LoadQueue.scala 314:36:@12914.6]
  assign _GEN_653 = initBits_4 ? 1'h0 : _GEN_652; // @[LoadQueue.scala 308:34:@12894.4]
  assign _GEN_654 = initBits_4 ? addrQ_4 : _GEN_651; // @[LoadQueue.scala 308:34:@12894.4]
  assign _T_31711 = inputPriorityPorts_0_5 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@12938.6]
  assign _T_31712 = inputPriorityPorts_1_5 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@12939.6]
  assign _T_31713 = inputPriorityPorts_2_5 & io_loadAddrEnable_2; // @[LoadQueue.scala 313:47:@12940.6]
  assign _T_31714 = inputPriorityPorts_3_5 & io_loadAddrEnable_3; // @[LoadQueue.scala 313:47:@12941.6]
  assign _T_31715 = inputPriorityPorts_4_5 & io_loadAddrEnable_4; // @[LoadQueue.scala 313:47:@12942.6]
  assign _T_31729 = _T_31711 | _T_31712; // @[LoadQueue.scala 314:26:@12950.6]
  assign _T_31730 = _T_31729 | _T_31713; // @[LoadQueue.scala 314:26:@12951.6]
  assign _T_31731 = _T_31730 | _T_31714; // @[LoadQueue.scala 314:26:@12952.6]
  assign _T_31732 = _T_31731 | _T_31715; // @[LoadQueue.scala 314:26:@12953.6]
  assign _T_31736 = {_T_31715,_T_31714,_T_31713,_T_31712,_T_31711}; // @[OneHot.scala 18:45:@12958.8]
  assign _T_31737 = _T_31736[4]; // @[OneHot.scala 26:18:@12959.8]
  assign _T_31738 = _T_31736[3:0]; // @[OneHot.scala 27:18:@12960.8]
  assign _GEN_819 = {{3'd0}, _T_31737}; // @[OneHot.scala 28:28:@12962.8]
  assign _T_31741 = _GEN_819 | _T_31738; // @[OneHot.scala 28:28:@12962.8]
  assign _T_31742 = _T_31741[3:2]; // @[OneHot.scala 26:18:@12963.8]
  assign _T_31743 = _T_31741[1:0]; // @[OneHot.scala 27:18:@12964.8]
  assign _T_31745 = _T_31742 != 2'h0; // @[OneHot.scala 28:14:@12965.8]
  assign _T_31746 = _T_31742 | _T_31743; // @[OneHot.scala 28:28:@12966.8]
  assign _T_31747 = _T_31746[1]; // @[CircuitMath.scala 30:8:@12967.8]
  assign _T_31749 = {_T_31737,_T_31745,_T_31747}; // @[Cat.scala 30:58:@12969.8]
  assign _GEN_656 = 3'h1 == _T_31749 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@12970.8]
  assign _GEN_657 = 3'h2 == _T_31749 ? io_addrFromLoadPorts_2 : _GEN_656; // @[LoadQueue.scala 315:29:@12970.8]
  assign _GEN_658 = 3'h3 == _T_31749 ? io_addrFromLoadPorts_3 : _GEN_657; // @[LoadQueue.scala 315:29:@12970.8]
  assign _GEN_659 = 3'h4 == _T_31749 ? io_addrFromLoadPorts_4 : _GEN_658; // @[LoadQueue.scala 315:29:@12970.8]
  assign _GEN_660 = _T_31732 ? _GEN_659 : addrQ_5; // @[LoadQueue.scala 314:36:@12954.6]
  assign _GEN_661 = _T_31732 ? 1'h1 : addrKnown_5; // @[LoadQueue.scala 314:36:@12954.6]
  assign _GEN_662 = initBits_5 ? 1'h0 : _GEN_661; // @[LoadQueue.scala 308:34:@12934.4]
  assign _GEN_663 = initBits_5 ? addrQ_5 : _GEN_660; // @[LoadQueue.scala 308:34:@12934.4]
  assign _T_31753 = inputPriorityPorts_0_6 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@12978.6]
  assign _T_31754 = inputPriorityPorts_1_6 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@12979.6]
  assign _T_31755 = inputPriorityPorts_2_6 & io_loadAddrEnable_2; // @[LoadQueue.scala 313:47:@12980.6]
  assign _T_31756 = inputPriorityPorts_3_6 & io_loadAddrEnable_3; // @[LoadQueue.scala 313:47:@12981.6]
  assign _T_31757 = inputPriorityPorts_4_6 & io_loadAddrEnable_4; // @[LoadQueue.scala 313:47:@12982.6]
  assign _T_31771 = _T_31753 | _T_31754; // @[LoadQueue.scala 314:26:@12990.6]
  assign _T_31772 = _T_31771 | _T_31755; // @[LoadQueue.scala 314:26:@12991.6]
  assign _T_31773 = _T_31772 | _T_31756; // @[LoadQueue.scala 314:26:@12992.6]
  assign _T_31774 = _T_31773 | _T_31757; // @[LoadQueue.scala 314:26:@12993.6]
  assign _T_31778 = {_T_31757,_T_31756,_T_31755,_T_31754,_T_31753}; // @[OneHot.scala 18:45:@12998.8]
  assign _T_31779 = _T_31778[4]; // @[OneHot.scala 26:18:@12999.8]
  assign _T_31780 = _T_31778[3:0]; // @[OneHot.scala 27:18:@13000.8]
  assign _GEN_820 = {{3'd0}, _T_31779}; // @[OneHot.scala 28:28:@13002.8]
  assign _T_31783 = _GEN_820 | _T_31780; // @[OneHot.scala 28:28:@13002.8]
  assign _T_31784 = _T_31783[3:2]; // @[OneHot.scala 26:18:@13003.8]
  assign _T_31785 = _T_31783[1:0]; // @[OneHot.scala 27:18:@13004.8]
  assign _T_31787 = _T_31784 != 2'h0; // @[OneHot.scala 28:14:@13005.8]
  assign _T_31788 = _T_31784 | _T_31785; // @[OneHot.scala 28:28:@13006.8]
  assign _T_31789 = _T_31788[1]; // @[CircuitMath.scala 30:8:@13007.8]
  assign _T_31791 = {_T_31779,_T_31787,_T_31789}; // @[Cat.scala 30:58:@13009.8]
  assign _GEN_665 = 3'h1 == _T_31791 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@13010.8]
  assign _GEN_666 = 3'h2 == _T_31791 ? io_addrFromLoadPorts_2 : _GEN_665; // @[LoadQueue.scala 315:29:@13010.8]
  assign _GEN_667 = 3'h3 == _T_31791 ? io_addrFromLoadPorts_3 : _GEN_666; // @[LoadQueue.scala 315:29:@13010.8]
  assign _GEN_668 = 3'h4 == _T_31791 ? io_addrFromLoadPorts_4 : _GEN_667; // @[LoadQueue.scala 315:29:@13010.8]
  assign _GEN_669 = _T_31774 ? _GEN_668 : addrQ_6; // @[LoadQueue.scala 314:36:@12994.6]
  assign _GEN_670 = _T_31774 ? 1'h1 : addrKnown_6; // @[LoadQueue.scala 314:36:@12994.6]
  assign _GEN_671 = initBits_6 ? 1'h0 : _GEN_670; // @[LoadQueue.scala 308:34:@12974.4]
  assign _GEN_672 = initBits_6 ? addrQ_6 : _GEN_669; // @[LoadQueue.scala 308:34:@12974.4]
  assign _T_31795 = inputPriorityPorts_0_7 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@13018.6]
  assign _T_31796 = inputPriorityPorts_1_7 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@13019.6]
  assign _T_31797 = inputPriorityPorts_2_7 & io_loadAddrEnable_2; // @[LoadQueue.scala 313:47:@13020.6]
  assign _T_31798 = inputPriorityPorts_3_7 & io_loadAddrEnable_3; // @[LoadQueue.scala 313:47:@13021.6]
  assign _T_31799 = inputPriorityPorts_4_7 & io_loadAddrEnable_4; // @[LoadQueue.scala 313:47:@13022.6]
  assign _T_31813 = _T_31795 | _T_31796; // @[LoadQueue.scala 314:26:@13030.6]
  assign _T_31814 = _T_31813 | _T_31797; // @[LoadQueue.scala 314:26:@13031.6]
  assign _T_31815 = _T_31814 | _T_31798; // @[LoadQueue.scala 314:26:@13032.6]
  assign _T_31816 = _T_31815 | _T_31799; // @[LoadQueue.scala 314:26:@13033.6]
  assign _T_31820 = {_T_31799,_T_31798,_T_31797,_T_31796,_T_31795}; // @[OneHot.scala 18:45:@13038.8]
  assign _T_31821 = _T_31820[4]; // @[OneHot.scala 26:18:@13039.8]
  assign _T_31822 = _T_31820[3:0]; // @[OneHot.scala 27:18:@13040.8]
  assign _GEN_821 = {{3'd0}, _T_31821}; // @[OneHot.scala 28:28:@13042.8]
  assign _T_31825 = _GEN_821 | _T_31822; // @[OneHot.scala 28:28:@13042.8]
  assign _T_31826 = _T_31825[3:2]; // @[OneHot.scala 26:18:@13043.8]
  assign _T_31827 = _T_31825[1:0]; // @[OneHot.scala 27:18:@13044.8]
  assign _T_31829 = _T_31826 != 2'h0; // @[OneHot.scala 28:14:@13045.8]
  assign _T_31830 = _T_31826 | _T_31827; // @[OneHot.scala 28:28:@13046.8]
  assign _T_31831 = _T_31830[1]; // @[CircuitMath.scala 30:8:@13047.8]
  assign _T_31833 = {_T_31821,_T_31829,_T_31831}; // @[Cat.scala 30:58:@13049.8]
  assign _GEN_674 = 3'h1 == _T_31833 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@13050.8]
  assign _GEN_675 = 3'h2 == _T_31833 ? io_addrFromLoadPorts_2 : _GEN_674; // @[LoadQueue.scala 315:29:@13050.8]
  assign _GEN_676 = 3'h3 == _T_31833 ? io_addrFromLoadPorts_3 : _GEN_675; // @[LoadQueue.scala 315:29:@13050.8]
  assign _GEN_677 = 3'h4 == _T_31833 ? io_addrFromLoadPorts_4 : _GEN_676; // @[LoadQueue.scala 315:29:@13050.8]
  assign _GEN_678 = _T_31816 ? _GEN_677 : addrQ_7; // @[LoadQueue.scala 314:36:@13034.6]
  assign _GEN_679 = _T_31816 ? 1'h1 : addrKnown_7; // @[LoadQueue.scala 314:36:@13034.6]
  assign _GEN_680 = initBits_7 ? 1'h0 : _GEN_679; // @[LoadQueue.scala 308:34:@13014.4]
  assign _GEN_681 = initBits_7 ? addrQ_7 : _GEN_678; // @[LoadQueue.scala 308:34:@13014.4]
  assign _T_31849 = outputPriorityPorts_0_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@13055.4]
  assign _T_31851 = loadCompleted_0 == 1'h0; // @[LoadQueue.scala 327:34:@13056.4]
  assign _T_31852 = _T_31849 & _T_31851; // @[LoadQueue.scala 327:31:@13057.4]
  assign _T_31853 = _T_31852 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@13058.4]
  assign _T_31854 = outputPriorityPorts_1_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@13059.4]
  assign _T_31857 = _T_31854 & _T_31851; // @[LoadQueue.scala 327:31:@13061.4]
  assign _T_31858 = _T_31857 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@13062.4]
  assign _T_31859 = outputPriorityPorts_2_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@13063.4]
  assign _T_31862 = _T_31859 & _T_31851; // @[LoadQueue.scala 327:31:@13065.4]
  assign _T_31863 = _T_31862 & io_loadPorts_2_ready; // @[LoadQueue.scala 327:63:@13066.4]
  assign _T_31864 = outputPriorityPorts_3_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@13067.4]
  assign _T_31867 = _T_31864 & _T_31851; // @[LoadQueue.scala 327:31:@13069.4]
  assign _T_31868 = _T_31867 & io_loadPorts_3_ready; // @[LoadQueue.scala 327:63:@13070.4]
  assign _T_31869 = outputPriorityPorts_4_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@13071.4]
  assign _T_31872 = _T_31869 & _T_31851; // @[LoadQueue.scala 327:31:@13073.4]
  assign _T_31873 = _T_31872 & io_loadPorts_4_ready; // @[LoadQueue.scala 327:63:@13074.4]
  assign _T_31887 = _T_31853 | _T_31858; // @[LoadQueue.scala 328:51:@13082.4]
  assign _T_31888 = _T_31887 | _T_31863; // @[LoadQueue.scala 328:51:@13083.4]
  assign _T_31889 = _T_31888 | _T_31868; // @[LoadQueue.scala 328:51:@13084.4]
  assign loadCompleting_0 = _T_31889 | _T_31873; // @[LoadQueue.scala 328:51:@13085.4]
  assign _T_31891 = outputPriorityPorts_0_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@13087.4]
  assign _T_31893 = loadCompleted_1 == 1'h0; // @[LoadQueue.scala 327:34:@13088.4]
  assign _T_31894 = _T_31891 & _T_31893; // @[LoadQueue.scala 327:31:@13089.4]
  assign _T_31895 = _T_31894 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@13090.4]
  assign _T_31896 = outputPriorityPorts_1_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@13091.4]
  assign _T_31899 = _T_31896 & _T_31893; // @[LoadQueue.scala 327:31:@13093.4]
  assign _T_31900 = _T_31899 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@13094.4]
  assign _T_31901 = outputPriorityPorts_2_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@13095.4]
  assign _T_31904 = _T_31901 & _T_31893; // @[LoadQueue.scala 327:31:@13097.4]
  assign _T_31905 = _T_31904 & io_loadPorts_2_ready; // @[LoadQueue.scala 327:63:@13098.4]
  assign _T_31906 = outputPriorityPorts_3_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@13099.4]
  assign _T_31909 = _T_31906 & _T_31893; // @[LoadQueue.scala 327:31:@13101.4]
  assign _T_31910 = _T_31909 & io_loadPorts_3_ready; // @[LoadQueue.scala 327:63:@13102.4]
  assign _T_31911 = outputPriorityPorts_4_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@13103.4]
  assign _T_31914 = _T_31911 & _T_31893; // @[LoadQueue.scala 327:31:@13105.4]
  assign _T_31915 = _T_31914 & io_loadPorts_4_ready; // @[LoadQueue.scala 327:63:@13106.4]
  assign _T_31929 = _T_31895 | _T_31900; // @[LoadQueue.scala 328:51:@13114.4]
  assign _T_31930 = _T_31929 | _T_31905; // @[LoadQueue.scala 328:51:@13115.4]
  assign _T_31931 = _T_31930 | _T_31910; // @[LoadQueue.scala 328:51:@13116.4]
  assign loadCompleting_1 = _T_31931 | _T_31915; // @[LoadQueue.scala 328:51:@13117.4]
  assign _T_31933 = outputPriorityPorts_0_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@13119.4]
  assign _T_31935 = loadCompleted_2 == 1'h0; // @[LoadQueue.scala 327:34:@13120.4]
  assign _T_31936 = _T_31933 & _T_31935; // @[LoadQueue.scala 327:31:@13121.4]
  assign _T_31937 = _T_31936 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@13122.4]
  assign _T_31938 = outputPriorityPorts_1_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@13123.4]
  assign _T_31941 = _T_31938 & _T_31935; // @[LoadQueue.scala 327:31:@13125.4]
  assign _T_31942 = _T_31941 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@13126.4]
  assign _T_31943 = outputPriorityPorts_2_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@13127.4]
  assign _T_31946 = _T_31943 & _T_31935; // @[LoadQueue.scala 327:31:@13129.4]
  assign _T_31947 = _T_31946 & io_loadPorts_2_ready; // @[LoadQueue.scala 327:63:@13130.4]
  assign _T_31948 = outputPriorityPorts_3_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@13131.4]
  assign _T_31951 = _T_31948 & _T_31935; // @[LoadQueue.scala 327:31:@13133.4]
  assign _T_31952 = _T_31951 & io_loadPorts_3_ready; // @[LoadQueue.scala 327:63:@13134.4]
  assign _T_31953 = outputPriorityPorts_4_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@13135.4]
  assign _T_31956 = _T_31953 & _T_31935; // @[LoadQueue.scala 327:31:@13137.4]
  assign _T_31957 = _T_31956 & io_loadPorts_4_ready; // @[LoadQueue.scala 327:63:@13138.4]
  assign _T_31971 = _T_31937 | _T_31942; // @[LoadQueue.scala 328:51:@13146.4]
  assign _T_31972 = _T_31971 | _T_31947; // @[LoadQueue.scala 328:51:@13147.4]
  assign _T_31973 = _T_31972 | _T_31952; // @[LoadQueue.scala 328:51:@13148.4]
  assign loadCompleting_2 = _T_31973 | _T_31957; // @[LoadQueue.scala 328:51:@13149.4]
  assign _T_31975 = outputPriorityPorts_0_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@13151.4]
  assign _T_31977 = loadCompleted_3 == 1'h0; // @[LoadQueue.scala 327:34:@13152.4]
  assign _T_31978 = _T_31975 & _T_31977; // @[LoadQueue.scala 327:31:@13153.4]
  assign _T_31979 = _T_31978 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@13154.4]
  assign _T_31980 = outputPriorityPorts_1_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@13155.4]
  assign _T_31983 = _T_31980 & _T_31977; // @[LoadQueue.scala 327:31:@13157.4]
  assign _T_31984 = _T_31983 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@13158.4]
  assign _T_31985 = outputPriorityPorts_2_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@13159.4]
  assign _T_31988 = _T_31985 & _T_31977; // @[LoadQueue.scala 327:31:@13161.4]
  assign _T_31989 = _T_31988 & io_loadPorts_2_ready; // @[LoadQueue.scala 327:63:@13162.4]
  assign _T_31990 = outputPriorityPorts_3_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@13163.4]
  assign _T_31993 = _T_31990 & _T_31977; // @[LoadQueue.scala 327:31:@13165.4]
  assign _T_31994 = _T_31993 & io_loadPorts_3_ready; // @[LoadQueue.scala 327:63:@13166.4]
  assign _T_31995 = outputPriorityPorts_4_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@13167.4]
  assign _T_31998 = _T_31995 & _T_31977; // @[LoadQueue.scala 327:31:@13169.4]
  assign _T_31999 = _T_31998 & io_loadPorts_4_ready; // @[LoadQueue.scala 327:63:@13170.4]
  assign _T_32013 = _T_31979 | _T_31984; // @[LoadQueue.scala 328:51:@13178.4]
  assign _T_32014 = _T_32013 | _T_31989; // @[LoadQueue.scala 328:51:@13179.4]
  assign _T_32015 = _T_32014 | _T_31994; // @[LoadQueue.scala 328:51:@13180.4]
  assign loadCompleting_3 = _T_32015 | _T_31999; // @[LoadQueue.scala 328:51:@13181.4]
  assign _T_32017 = outputPriorityPorts_0_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@13183.4]
  assign _T_32019 = loadCompleted_4 == 1'h0; // @[LoadQueue.scala 327:34:@13184.4]
  assign _T_32020 = _T_32017 & _T_32019; // @[LoadQueue.scala 327:31:@13185.4]
  assign _T_32021 = _T_32020 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@13186.4]
  assign _T_32022 = outputPriorityPorts_1_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@13187.4]
  assign _T_32025 = _T_32022 & _T_32019; // @[LoadQueue.scala 327:31:@13189.4]
  assign _T_32026 = _T_32025 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@13190.4]
  assign _T_32027 = outputPriorityPorts_2_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@13191.4]
  assign _T_32030 = _T_32027 & _T_32019; // @[LoadQueue.scala 327:31:@13193.4]
  assign _T_32031 = _T_32030 & io_loadPorts_2_ready; // @[LoadQueue.scala 327:63:@13194.4]
  assign _T_32032 = outputPriorityPorts_3_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@13195.4]
  assign _T_32035 = _T_32032 & _T_32019; // @[LoadQueue.scala 327:31:@13197.4]
  assign _T_32036 = _T_32035 & io_loadPorts_3_ready; // @[LoadQueue.scala 327:63:@13198.4]
  assign _T_32037 = outputPriorityPorts_4_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@13199.4]
  assign _T_32040 = _T_32037 & _T_32019; // @[LoadQueue.scala 327:31:@13201.4]
  assign _T_32041 = _T_32040 & io_loadPorts_4_ready; // @[LoadQueue.scala 327:63:@13202.4]
  assign _T_32055 = _T_32021 | _T_32026; // @[LoadQueue.scala 328:51:@13210.4]
  assign _T_32056 = _T_32055 | _T_32031; // @[LoadQueue.scala 328:51:@13211.4]
  assign _T_32057 = _T_32056 | _T_32036; // @[LoadQueue.scala 328:51:@13212.4]
  assign loadCompleting_4 = _T_32057 | _T_32041; // @[LoadQueue.scala 328:51:@13213.4]
  assign _T_32059 = outputPriorityPorts_0_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@13215.4]
  assign _T_32061 = loadCompleted_5 == 1'h0; // @[LoadQueue.scala 327:34:@13216.4]
  assign _T_32062 = _T_32059 & _T_32061; // @[LoadQueue.scala 327:31:@13217.4]
  assign _T_32063 = _T_32062 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@13218.4]
  assign _T_32064 = outputPriorityPorts_1_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@13219.4]
  assign _T_32067 = _T_32064 & _T_32061; // @[LoadQueue.scala 327:31:@13221.4]
  assign _T_32068 = _T_32067 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@13222.4]
  assign _T_32069 = outputPriorityPorts_2_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@13223.4]
  assign _T_32072 = _T_32069 & _T_32061; // @[LoadQueue.scala 327:31:@13225.4]
  assign _T_32073 = _T_32072 & io_loadPorts_2_ready; // @[LoadQueue.scala 327:63:@13226.4]
  assign _T_32074 = outputPriorityPorts_3_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@13227.4]
  assign _T_32077 = _T_32074 & _T_32061; // @[LoadQueue.scala 327:31:@13229.4]
  assign _T_32078 = _T_32077 & io_loadPorts_3_ready; // @[LoadQueue.scala 327:63:@13230.4]
  assign _T_32079 = outputPriorityPorts_4_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@13231.4]
  assign _T_32082 = _T_32079 & _T_32061; // @[LoadQueue.scala 327:31:@13233.4]
  assign _T_32083 = _T_32082 & io_loadPorts_4_ready; // @[LoadQueue.scala 327:63:@13234.4]
  assign _T_32097 = _T_32063 | _T_32068; // @[LoadQueue.scala 328:51:@13242.4]
  assign _T_32098 = _T_32097 | _T_32073; // @[LoadQueue.scala 328:51:@13243.4]
  assign _T_32099 = _T_32098 | _T_32078; // @[LoadQueue.scala 328:51:@13244.4]
  assign loadCompleting_5 = _T_32099 | _T_32083; // @[LoadQueue.scala 328:51:@13245.4]
  assign _T_32101 = outputPriorityPorts_0_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@13247.4]
  assign _T_32103 = loadCompleted_6 == 1'h0; // @[LoadQueue.scala 327:34:@13248.4]
  assign _T_32104 = _T_32101 & _T_32103; // @[LoadQueue.scala 327:31:@13249.4]
  assign _T_32105 = _T_32104 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@13250.4]
  assign _T_32106 = outputPriorityPorts_1_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@13251.4]
  assign _T_32109 = _T_32106 & _T_32103; // @[LoadQueue.scala 327:31:@13253.4]
  assign _T_32110 = _T_32109 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@13254.4]
  assign _T_32111 = outputPriorityPorts_2_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@13255.4]
  assign _T_32114 = _T_32111 & _T_32103; // @[LoadQueue.scala 327:31:@13257.4]
  assign _T_32115 = _T_32114 & io_loadPorts_2_ready; // @[LoadQueue.scala 327:63:@13258.4]
  assign _T_32116 = outputPriorityPorts_3_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@13259.4]
  assign _T_32119 = _T_32116 & _T_32103; // @[LoadQueue.scala 327:31:@13261.4]
  assign _T_32120 = _T_32119 & io_loadPorts_3_ready; // @[LoadQueue.scala 327:63:@13262.4]
  assign _T_32121 = outputPriorityPorts_4_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@13263.4]
  assign _T_32124 = _T_32121 & _T_32103; // @[LoadQueue.scala 327:31:@13265.4]
  assign _T_32125 = _T_32124 & io_loadPorts_4_ready; // @[LoadQueue.scala 327:63:@13266.4]
  assign _T_32139 = _T_32105 | _T_32110; // @[LoadQueue.scala 328:51:@13274.4]
  assign _T_32140 = _T_32139 | _T_32115; // @[LoadQueue.scala 328:51:@13275.4]
  assign _T_32141 = _T_32140 | _T_32120; // @[LoadQueue.scala 328:51:@13276.4]
  assign loadCompleting_6 = _T_32141 | _T_32125; // @[LoadQueue.scala 328:51:@13277.4]
  assign _T_32143 = outputPriorityPorts_0_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@13279.4]
  assign _T_32145 = loadCompleted_7 == 1'h0; // @[LoadQueue.scala 327:34:@13280.4]
  assign _T_32146 = _T_32143 & _T_32145; // @[LoadQueue.scala 327:31:@13281.4]
  assign _T_32147 = _T_32146 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@13282.4]
  assign _T_32148 = outputPriorityPorts_1_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@13283.4]
  assign _T_32151 = _T_32148 & _T_32145; // @[LoadQueue.scala 327:31:@13285.4]
  assign _T_32152 = _T_32151 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@13286.4]
  assign _T_32153 = outputPriorityPorts_2_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@13287.4]
  assign _T_32156 = _T_32153 & _T_32145; // @[LoadQueue.scala 327:31:@13289.4]
  assign _T_32157 = _T_32156 & io_loadPorts_2_ready; // @[LoadQueue.scala 327:63:@13290.4]
  assign _T_32158 = outputPriorityPorts_3_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@13291.4]
  assign _T_32161 = _T_32158 & _T_32145; // @[LoadQueue.scala 327:31:@13293.4]
  assign _T_32162 = _T_32161 & io_loadPorts_3_ready; // @[LoadQueue.scala 327:63:@13294.4]
  assign _T_32163 = outputPriorityPorts_4_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@13295.4]
  assign _T_32166 = _T_32163 & _T_32145; // @[LoadQueue.scala 327:31:@13297.4]
  assign _T_32167 = _T_32166 & io_loadPorts_4_ready; // @[LoadQueue.scala 327:63:@13298.4]
  assign _T_32181 = _T_32147 | _T_32152; // @[LoadQueue.scala 328:51:@13306.4]
  assign _T_32182 = _T_32181 | _T_32157; // @[LoadQueue.scala 328:51:@13307.4]
  assign _T_32183 = _T_32182 | _T_32162; // @[LoadQueue.scala 328:51:@13308.4]
  assign loadCompleting_7 = _T_32183 | _T_32167; // @[LoadQueue.scala 328:51:@13309.4]
  assign _GEN_682 = loadCompleting_0 ? 1'h1 : loadCompleted_0; // @[LoadQueue.scala 337:46:@13315.6]
  assign _GEN_683 = initBits_0 ? 1'h0 : _GEN_682; // @[LoadQueue.scala 335:34:@13311.4]
  assign _GEN_684 = loadCompleting_1 ? 1'h1 : loadCompleted_1; // @[LoadQueue.scala 337:46:@13322.6]
  assign _GEN_685 = initBits_1 ? 1'h0 : _GEN_684; // @[LoadQueue.scala 335:34:@13318.4]
  assign _GEN_686 = loadCompleting_2 ? 1'h1 : loadCompleted_2; // @[LoadQueue.scala 337:46:@13329.6]
  assign _GEN_687 = initBits_2 ? 1'h0 : _GEN_686; // @[LoadQueue.scala 335:34:@13325.4]
  assign _GEN_688 = loadCompleting_3 ? 1'h1 : loadCompleted_3; // @[LoadQueue.scala 337:46:@13336.6]
  assign _GEN_689 = initBits_3 ? 1'h0 : _GEN_688; // @[LoadQueue.scala 335:34:@13332.4]
  assign _GEN_690 = loadCompleting_4 ? 1'h1 : loadCompleted_4; // @[LoadQueue.scala 337:46:@13343.6]
  assign _GEN_691 = initBits_4 ? 1'h0 : _GEN_690; // @[LoadQueue.scala 335:34:@13339.4]
  assign _GEN_692 = loadCompleting_5 ? 1'h1 : loadCompleted_5; // @[LoadQueue.scala 337:46:@13350.6]
  assign _GEN_693 = initBits_5 ? 1'h0 : _GEN_692; // @[LoadQueue.scala 335:34:@13346.4]
  assign _GEN_694 = loadCompleting_6 ? 1'h1 : loadCompleted_6; // @[LoadQueue.scala 337:46:@13357.6]
  assign _GEN_695 = initBits_6 ? 1'h0 : _GEN_694; // @[LoadQueue.scala 335:34:@13353.4]
  assign _GEN_696 = loadCompleting_7 ? 1'h1 : loadCompleted_7; // @[LoadQueue.scala 337:46:@13364.6]
  assign _GEN_697 = initBits_7 ? 1'h0 : _GEN_696; // @[LoadQueue.scala 335:34:@13360.4]
  assign _T_32249 = _T_31852 | _T_31894; // @[LoadQueue.scala 348:24:@13401.4]
  assign _T_32250 = _T_32249 | _T_31936; // @[LoadQueue.scala 348:24:@13402.4]
  assign _T_32251 = _T_32250 | _T_31978; // @[LoadQueue.scala 348:24:@13403.4]
  assign _T_32252 = _T_32251 | _T_32020; // @[LoadQueue.scala 348:24:@13404.4]
  assign _T_32253 = _T_32252 | _T_32062; // @[LoadQueue.scala 348:24:@13405.4]
  assign _T_32254 = _T_32253 | _T_32104; // @[LoadQueue.scala 348:24:@13406.4]
  assign _T_32255 = _T_32254 | _T_32146; // @[LoadQueue.scala 348:24:@13407.4]
  assign _T_32264 = _T_32104 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@13409.6]
  assign _T_32265 = _T_32062 ? 3'h5 : _T_32264; // @[Mux.scala 31:69:@13410.6]
  assign _T_32266 = _T_32020 ? 3'h4 : _T_32265; // @[Mux.scala 31:69:@13411.6]
  assign _T_32267 = _T_31978 ? 3'h3 : _T_32266; // @[Mux.scala 31:69:@13412.6]
  assign _T_32268 = _T_31936 ? 3'h2 : _T_32267; // @[Mux.scala 31:69:@13413.6]
  assign _T_32269 = _T_31894 ? 3'h1 : _T_32268; // @[Mux.scala 31:69:@13414.6]
  assign _T_32270 = _T_31852 ? 3'h0 : _T_32269; // @[Mux.scala 31:69:@13415.6]
  assign _GEN_699 = 3'h1 == _T_32270 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@13416.6]
  assign _GEN_700 = 3'h2 == _T_32270 ? dataQ_2 : _GEN_699; // @[LoadQueue.scala 349:37:@13416.6]
  assign _GEN_701 = 3'h3 == _T_32270 ? dataQ_3 : _GEN_700; // @[LoadQueue.scala 349:37:@13416.6]
  assign _GEN_702 = 3'h4 == _T_32270 ? dataQ_4 : _GEN_701; // @[LoadQueue.scala 349:37:@13416.6]
  assign _GEN_703 = 3'h5 == _T_32270 ? dataQ_5 : _GEN_702; // @[LoadQueue.scala 349:37:@13416.6]
  assign _GEN_704 = 3'h6 == _T_32270 ? dataQ_6 : _GEN_703; // @[LoadQueue.scala 349:37:@13416.6]
  assign _GEN_705 = 3'h7 == _T_32270 ? dataQ_7 : _GEN_704; // @[LoadQueue.scala 349:37:@13416.6]
  assign _T_32325 = _T_31857 | _T_31899; // @[LoadQueue.scala 348:24:@13457.4]
  assign _T_32326 = _T_32325 | _T_31941; // @[LoadQueue.scala 348:24:@13458.4]
  assign _T_32327 = _T_32326 | _T_31983; // @[LoadQueue.scala 348:24:@13459.4]
  assign _T_32328 = _T_32327 | _T_32025; // @[LoadQueue.scala 348:24:@13460.4]
  assign _T_32329 = _T_32328 | _T_32067; // @[LoadQueue.scala 348:24:@13461.4]
  assign _T_32330 = _T_32329 | _T_32109; // @[LoadQueue.scala 348:24:@13462.4]
  assign _T_32331 = _T_32330 | _T_32151; // @[LoadQueue.scala 348:24:@13463.4]
  assign _T_32340 = _T_32109 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@13465.6]
  assign _T_32341 = _T_32067 ? 3'h5 : _T_32340; // @[Mux.scala 31:69:@13466.6]
  assign _T_32342 = _T_32025 ? 3'h4 : _T_32341; // @[Mux.scala 31:69:@13467.6]
  assign _T_32343 = _T_31983 ? 3'h3 : _T_32342; // @[Mux.scala 31:69:@13468.6]
  assign _T_32344 = _T_31941 ? 3'h2 : _T_32343; // @[Mux.scala 31:69:@13469.6]
  assign _T_32345 = _T_31899 ? 3'h1 : _T_32344; // @[Mux.scala 31:69:@13470.6]
  assign _T_32346 = _T_31857 ? 3'h0 : _T_32345; // @[Mux.scala 31:69:@13471.6]
  assign _GEN_709 = 3'h1 == _T_32346 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@13472.6]
  assign _GEN_710 = 3'h2 == _T_32346 ? dataQ_2 : _GEN_709; // @[LoadQueue.scala 349:37:@13472.6]
  assign _GEN_711 = 3'h3 == _T_32346 ? dataQ_3 : _GEN_710; // @[LoadQueue.scala 349:37:@13472.6]
  assign _GEN_712 = 3'h4 == _T_32346 ? dataQ_4 : _GEN_711; // @[LoadQueue.scala 349:37:@13472.6]
  assign _GEN_713 = 3'h5 == _T_32346 ? dataQ_5 : _GEN_712; // @[LoadQueue.scala 349:37:@13472.6]
  assign _GEN_714 = 3'h6 == _T_32346 ? dataQ_6 : _GEN_713; // @[LoadQueue.scala 349:37:@13472.6]
  assign _GEN_715 = 3'h7 == _T_32346 ? dataQ_7 : _GEN_714; // @[LoadQueue.scala 349:37:@13472.6]
  assign _T_32401 = _T_31862 | _T_31904; // @[LoadQueue.scala 348:24:@13513.4]
  assign _T_32402 = _T_32401 | _T_31946; // @[LoadQueue.scala 348:24:@13514.4]
  assign _T_32403 = _T_32402 | _T_31988; // @[LoadQueue.scala 348:24:@13515.4]
  assign _T_32404 = _T_32403 | _T_32030; // @[LoadQueue.scala 348:24:@13516.4]
  assign _T_32405 = _T_32404 | _T_32072; // @[LoadQueue.scala 348:24:@13517.4]
  assign _T_32406 = _T_32405 | _T_32114; // @[LoadQueue.scala 348:24:@13518.4]
  assign _T_32407 = _T_32406 | _T_32156; // @[LoadQueue.scala 348:24:@13519.4]
  assign _T_32416 = _T_32114 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@13521.6]
  assign _T_32417 = _T_32072 ? 3'h5 : _T_32416; // @[Mux.scala 31:69:@13522.6]
  assign _T_32418 = _T_32030 ? 3'h4 : _T_32417; // @[Mux.scala 31:69:@13523.6]
  assign _T_32419 = _T_31988 ? 3'h3 : _T_32418; // @[Mux.scala 31:69:@13524.6]
  assign _T_32420 = _T_31946 ? 3'h2 : _T_32419; // @[Mux.scala 31:69:@13525.6]
  assign _T_32421 = _T_31904 ? 3'h1 : _T_32420; // @[Mux.scala 31:69:@13526.6]
  assign _T_32422 = _T_31862 ? 3'h0 : _T_32421; // @[Mux.scala 31:69:@13527.6]
  assign _GEN_719 = 3'h1 == _T_32422 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@13528.6]
  assign _GEN_720 = 3'h2 == _T_32422 ? dataQ_2 : _GEN_719; // @[LoadQueue.scala 349:37:@13528.6]
  assign _GEN_721 = 3'h3 == _T_32422 ? dataQ_3 : _GEN_720; // @[LoadQueue.scala 349:37:@13528.6]
  assign _GEN_722 = 3'h4 == _T_32422 ? dataQ_4 : _GEN_721; // @[LoadQueue.scala 349:37:@13528.6]
  assign _GEN_723 = 3'h5 == _T_32422 ? dataQ_5 : _GEN_722; // @[LoadQueue.scala 349:37:@13528.6]
  assign _GEN_724 = 3'h6 == _T_32422 ? dataQ_6 : _GEN_723; // @[LoadQueue.scala 349:37:@13528.6]
  assign _GEN_725 = 3'h7 == _T_32422 ? dataQ_7 : _GEN_724; // @[LoadQueue.scala 349:37:@13528.6]
  assign _T_32477 = _T_31867 | _T_31909; // @[LoadQueue.scala 348:24:@13569.4]
  assign _T_32478 = _T_32477 | _T_31951; // @[LoadQueue.scala 348:24:@13570.4]
  assign _T_32479 = _T_32478 | _T_31993; // @[LoadQueue.scala 348:24:@13571.4]
  assign _T_32480 = _T_32479 | _T_32035; // @[LoadQueue.scala 348:24:@13572.4]
  assign _T_32481 = _T_32480 | _T_32077; // @[LoadQueue.scala 348:24:@13573.4]
  assign _T_32482 = _T_32481 | _T_32119; // @[LoadQueue.scala 348:24:@13574.4]
  assign _T_32483 = _T_32482 | _T_32161; // @[LoadQueue.scala 348:24:@13575.4]
  assign _T_32492 = _T_32119 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@13577.6]
  assign _T_32493 = _T_32077 ? 3'h5 : _T_32492; // @[Mux.scala 31:69:@13578.6]
  assign _T_32494 = _T_32035 ? 3'h4 : _T_32493; // @[Mux.scala 31:69:@13579.6]
  assign _T_32495 = _T_31993 ? 3'h3 : _T_32494; // @[Mux.scala 31:69:@13580.6]
  assign _T_32496 = _T_31951 ? 3'h2 : _T_32495; // @[Mux.scala 31:69:@13581.6]
  assign _T_32497 = _T_31909 ? 3'h1 : _T_32496; // @[Mux.scala 31:69:@13582.6]
  assign _T_32498 = _T_31867 ? 3'h0 : _T_32497; // @[Mux.scala 31:69:@13583.6]
  assign _GEN_729 = 3'h1 == _T_32498 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@13584.6]
  assign _GEN_730 = 3'h2 == _T_32498 ? dataQ_2 : _GEN_729; // @[LoadQueue.scala 349:37:@13584.6]
  assign _GEN_731 = 3'h3 == _T_32498 ? dataQ_3 : _GEN_730; // @[LoadQueue.scala 349:37:@13584.6]
  assign _GEN_732 = 3'h4 == _T_32498 ? dataQ_4 : _GEN_731; // @[LoadQueue.scala 349:37:@13584.6]
  assign _GEN_733 = 3'h5 == _T_32498 ? dataQ_5 : _GEN_732; // @[LoadQueue.scala 349:37:@13584.6]
  assign _GEN_734 = 3'h6 == _T_32498 ? dataQ_6 : _GEN_733; // @[LoadQueue.scala 349:37:@13584.6]
  assign _GEN_735 = 3'h7 == _T_32498 ? dataQ_7 : _GEN_734; // @[LoadQueue.scala 349:37:@13584.6]
  assign _T_32553 = _T_31872 | _T_31914; // @[LoadQueue.scala 348:24:@13625.4]
  assign _T_32554 = _T_32553 | _T_31956; // @[LoadQueue.scala 348:24:@13626.4]
  assign _T_32555 = _T_32554 | _T_31998; // @[LoadQueue.scala 348:24:@13627.4]
  assign _T_32556 = _T_32555 | _T_32040; // @[LoadQueue.scala 348:24:@13628.4]
  assign _T_32557 = _T_32556 | _T_32082; // @[LoadQueue.scala 348:24:@13629.4]
  assign _T_32558 = _T_32557 | _T_32124; // @[LoadQueue.scala 348:24:@13630.4]
  assign _T_32559 = _T_32558 | _T_32166; // @[LoadQueue.scala 348:24:@13631.4]
  assign _T_32568 = _T_32124 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@13633.6]
  assign _T_32569 = _T_32082 ? 3'h5 : _T_32568; // @[Mux.scala 31:69:@13634.6]
  assign _T_32570 = _T_32040 ? 3'h4 : _T_32569; // @[Mux.scala 31:69:@13635.6]
  assign _T_32571 = _T_31998 ? 3'h3 : _T_32570; // @[Mux.scala 31:69:@13636.6]
  assign _T_32572 = _T_31956 ? 3'h2 : _T_32571; // @[Mux.scala 31:69:@13637.6]
  assign _T_32573 = _T_31914 ? 3'h1 : _T_32572; // @[Mux.scala 31:69:@13638.6]
  assign _T_32574 = _T_31872 ? 3'h0 : _T_32573; // @[Mux.scala 31:69:@13639.6]
  assign _GEN_739 = 3'h1 == _T_32574 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@13640.6]
  assign _GEN_740 = 3'h2 == _T_32574 ? dataQ_2 : _GEN_739; // @[LoadQueue.scala 349:37:@13640.6]
  assign _GEN_741 = 3'h3 == _T_32574 ? dataQ_3 : _GEN_740; // @[LoadQueue.scala 349:37:@13640.6]
  assign _GEN_742 = 3'h4 == _T_32574 ? dataQ_4 : _GEN_741; // @[LoadQueue.scala 349:37:@13640.6]
  assign _GEN_743 = 3'h5 == _T_32574 ? dataQ_5 : _GEN_742; // @[LoadQueue.scala 349:37:@13640.6]
  assign _GEN_744 = 3'h6 == _T_32574 ? dataQ_6 : _GEN_743; // @[LoadQueue.scala 349:37:@13640.6]
  assign _GEN_745 = 3'h7 == _T_32574 ? dataQ_7 : _GEN_744; // @[LoadQueue.scala 349:37:@13640.6]
  assign _GEN_749 = 3'h1 == head ? loadCompleted_1 : loadCompleted_0; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_750 = 3'h2 == head ? loadCompleted_2 : _GEN_749; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_751 = 3'h3 == head ? loadCompleted_3 : _GEN_750; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_752 = 3'h4 == head ? loadCompleted_4 : _GEN_751; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_753 = 3'h5 == head ? loadCompleted_5 : _GEN_752; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_754 = 3'h6 == head ? loadCompleted_6 : _GEN_753; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_755 = 3'h7 == head ? loadCompleted_7 : _GEN_754; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_757 = 3'h1 == head ? loadCompleting_1 : loadCompleting_0; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_758 = 3'h2 == head ? loadCompleting_2 : _GEN_757; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_759 = 3'h3 == head ? loadCompleting_3 : _GEN_758; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_760 = 3'h4 == head ? loadCompleting_4 : _GEN_759; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_761 = 3'h5 == head ? loadCompleting_5 : _GEN_760; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_762 = 3'h6 == head ? loadCompleting_6 : _GEN_761; // @[LoadQueue.scala 363:29:@13647.4]
  assign _GEN_763 = 3'h7 == head ? loadCompleting_7 : _GEN_762; // @[LoadQueue.scala 363:29:@13647.4]
  assign _T_32585 = _GEN_755 | _GEN_763; // @[LoadQueue.scala 363:29:@13647.4]
  assign _T_32586 = head != tail; // @[LoadQueue.scala 363:63:@13648.4]
  assign _T_32588 = io_loadEmpty == 1'h0; // @[LoadQueue.scala 363:75:@13649.4]
  assign _T_32589 = _T_32586 | _T_32588; // @[LoadQueue.scala 363:72:@13650.4]
  assign _T_32590 = _T_32585 & _T_32589; // @[LoadQueue.scala 363:54:@13651.4]
  assign _T_32593 = head + 3'h1; // @[util.scala 10:8:@13653.6]
  assign _GEN_144 = _T_32593 % 4'h8; // @[util.scala 10:14:@13654.6]
  assign _T_32594 = _GEN_144[3:0]; // @[util.scala 10:14:@13654.6]
  assign _GEN_764 = _T_32590 ? _T_32594 : {{1'd0}, head}; // @[LoadQueue.scala 363:91:@13652.4]
  assign _T_32596 = tail + io_bbNumLoads; // @[util.scala 10:8:@13658.6]
  assign _GEN_145 = _T_32596 % 4'h8; // @[util.scala 10:14:@13659.6]
  assign _T_32597 = _GEN_145[3:0]; // @[util.scala 10:14:@13659.6]
  assign _GEN_765 = io_bbStart ? _T_32597 : {{1'd0}, tail}; // @[LoadQueue.scala 367:20:@13657.4]
  assign _T_32599 = allocatedEntries_0 == 1'h0; // @[LoadQueue.scala 371:82:@13662.4]
  assign _T_32600 = loadCompleted_0 | _T_32599; // @[LoadQueue.scala 371:79:@13663.4]
  assign _T_32602 = allocatedEntries_1 == 1'h0; // @[LoadQueue.scala 371:82:@13664.4]
  assign _T_32603 = loadCompleted_1 | _T_32602; // @[LoadQueue.scala 371:79:@13665.4]
  assign _T_32605 = allocatedEntries_2 == 1'h0; // @[LoadQueue.scala 371:82:@13666.4]
  assign _T_32606 = loadCompleted_2 | _T_32605; // @[LoadQueue.scala 371:79:@13667.4]
  assign _T_32608 = allocatedEntries_3 == 1'h0; // @[LoadQueue.scala 371:82:@13668.4]
  assign _T_32609 = loadCompleted_3 | _T_32608; // @[LoadQueue.scala 371:79:@13669.4]
  assign _T_32611 = allocatedEntries_4 == 1'h0; // @[LoadQueue.scala 371:82:@13670.4]
  assign _T_32612 = loadCompleted_4 | _T_32611; // @[LoadQueue.scala 371:79:@13671.4]
  assign _T_32614 = allocatedEntries_5 == 1'h0; // @[LoadQueue.scala 371:82:@13672.4]
  assign _T_32615 = loadCompleted_5 | _T_32614; // @[LoadQueue.scala 371:79:@13673.4]
  assign _T_32617 = allocatedEntries_6 == 1'h0; // @[LoadQueue.scala 371:82:@13674.4]
  assign _T_32618 = loadCompleted_6 | _T_32617; // @[LoadQueue.scala 371:79:@13675.4]
  assign _T_32620 = allocatedEntries_7 == 1'h0; // @[LoadQueue.scala 371:82:@13676.4]
  assign _T_32621 = loadCompleted_7 | _T_32620; // @[LoadQueue.scala 371:79:@13677.4]
  assign _T_32638 = _T_32600 & _T_32603; // @[LoadQueue.scala 371:96:@13688.4]
  assign _T_32639 = _T_32638 & _T_32606; // @[LoadQueue.scala 371:96:@13689.4]
  assign _T_32640 = _T_32639 & _T_32609; // @[LoadQueue.scala 371:96:@13690.4]
  assign _T_32641 = _T_32640 & _T_32612; // @[LoadQueue.scala 371:96:@13691.4]
  assign _T_32642 = _T_32641 & _T_32615; // @[LoadQueue.scala 371:96:@13692.4]
  assign _T_32643 = _T_32642 & _T_32618; // @[LoadQueue.scala 371:96:@13693.4]
  assign io_loadTail = tail; // @[LoadQueue.scala 380:15:@13697.4]
  assign io_loadHead = head; // @[LoadQueue.scala 379:15:@13696.4]
  assign io_loadEmpty = _T_32643 & _T_32621; // @[LoadQueue.scala 371:16:@13695.4]
  assign io_loadAddrDone_0 = addrKnown_0; // @[LoadQueue.scala 382:19:@13706.4]
  assign io_loadAddrDone_1 = addrKnown_1; // @[LoadQueue.scala 382:19:@13707.4]
  assign io_loadAddrDone_2 = addrKnown_2; // @[LoadQueue.scala 382:19:@13708.4]
  assign io_loadAddrDone_3 = addrKnown_3; // @[LoadQueue.scala 382:19:@13709.4]
  assign io_loadAddrDone_4 = addrKnown_4; // @[LoadQueue.scala 382:19:@13710.4]
  assign io_loadAddrDone_5 = addrKnown_5; // @[LoadQueue.scala 382:19:@13711.4]
  assign io_loadAddrDone_6 = addrKnown_6; // @[LoadQueue.scala 382:19:@13712.4]
  assign io_loadAddrDone_7 = addrKnown_7; // @[LoadQueue.scala 382:19:@13713.4]
  assign io_loadDataDone_0 = dataKnown_0; // @[LoadQueue.scala 383:19:@13714.4]
  assign io_loadDataDone_1 = dataKnown_1; // @[LoadQueue.scala 383:19:@13715.4]
  assign io_loadDataDone_2 = dataKnown_2; // @[LoadQueue.scala 383:19:@13716.4]
  assign io_loadDataDone_3 = dataKnown_3; // @[LoadQueue.scala 383:19:@13717.4]
  assign io_loadDataDone_4 = dataKnown_4; // @[LoadQueue.scala 383:19:@13718.4]
  assign io_loadDataDone_5 = dataKnown_5; // @[LoadQueue.scala 383:19:@13719.4]
  assign io_loadDataDone_6 = dataKnown_6; // @[LoadQueue.scala 383:19:@13720.4]
  assign io_loadDataDone_7 = dataKnown_7; // @[LoadQueue.scala 383:19:@13721.4]
  assign io_loadAddrQueue_0 = addrQ_0; // @[LoadQueue.scala 381:20:@13698.4]
  assign io_loadAddrQueue_1 = addrQ_1; // @[LoadQueue.scala 381:20:@13699.4]
  assign io_loadAddrQueue_2 = addrQ_2; // @[LoadQueue.scala 381:20:@13700.4]
  assign io_loadAddrQueue_3 = addrQ_3; // @[LoadQueue.scala 381:20:@13701.4]
  assign io_loadAddrQueue_4 = addrQ_4; // @[LoadQueue.scala 381:20:@13702.4]
  assign io_loadAddrQueue_5 = addrQ_5; // @[LoadQueue.scala 381:20:@13703.4]
  assign io_loadAddrQueue_6 = addrQ_6; // @[LoadQueue.scala 381:20:@13704.4]
  assign io_loadAddrQueue_7 = addrQ_7; // @[LoadQueue.scala 381:20:@13705.4]
  assign io_loadPorts_0_valid = _T_32254 | _T_32146; // @[LoadQueue.scala 350:38:@13417.6 LoadQueue.scala 353:38:@13421.6]
  assign io_loadPorts_0_bits = _T_32255 ? _GEN_705 : 32'h0; // @[LoadQueue.scala 349:37:@13416.6 LoadQueue.scala 352:37:@13420.6]
  assign io_loadPorts_1_valid = _T_32330 | _T_32151; // @[LoadQueue.scala 350:38:@13473.6 LoadQueue.scala 353:38:@13477.6]
  assign io_loadPorts_1_bits = _T_32331 ? _GEN_715 : 32'h0; // @[LoadQueue.scala 349:37:@13472.6 LoadQueue.scala 352:37:@13476.6]
  assign io_loadPorts_2_valid = _T_32406 | _T_32156; // @[LoadQueue.scala 350:38:@13529.6 LoadQueue.scala 353:38:@13533.6]
  assign io_loadPorts_2_bits = _T_32407 ? _GEN_725 : 32'h0; // @[LoadQueue.scala 349:37:@13528.6 LoadQueue.scala 352:37:@13532.6]
  assign io_loadPorts_3_valid = _T_32482 | _T_32161; // @[LoadQueue.scala 350:38:@13585.6 LoadQueue.scala 353:38:@13589.6]
  assign io_loadPorts_3_bits = _T_32483 ? _GEN_735 : 32'h0; // @[LoadQueue.scala 349:37:@13584.6 LoadQueue.scala 352:37:@13588.6]
  assign io_loadPorts_4_valid = _T_32558 | _T_32166; // @[LoadQueue.scala 350:38:@13641.6 LoadQueue.scala 353:38:@13645.6]
  assign io_loadPorts_4_bits = _T_32559 ? _GEN_745 : 32'h0; // @[LoadQueue.scala 349:37:@13640.6 LoadQueue.scala 352:37:@13644.6]
  assign io_loadAddrToMem = _T_25226 ? _GEN_575 : 32'h0; // @[LoadQueue.scala 248:24:@9219.6 LoadQueue.scala 251:24:@9223.6]
  assign io_loadEnableToMem = _T_25225 | loadRequest_7; // @[LoadQueue.scala 246:22:@9202.4 LoadQueue.scala 249:26:@9220.6 LoadQueue.scala 252:26:@9224.6]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  portQ_0 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  portQ_1 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  portQ_2 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  portQ_3 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  portQ_4 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  portQ_5 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  portQ_6 = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  portQ_7 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  addrQ_0 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  addrQ_1 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  addrQ_2 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  addrQ_3 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  addrQ_4 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  addrQ_5 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  addrQ_6 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  addrQ_7 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  dataQ_0 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  dataQ_1 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  dataQ_2 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  dataQ_3 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  dataQ_4 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  dataQ_5 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  dataQ_6 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  dataQ_7 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrKnown_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrKnown_1 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrKnown_2 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrKnown_3 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrKnown_4 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrKnown_5 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrKnown_6 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrKnown_7 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  dataKnown_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  dataKnown_1 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  dataKnown_2 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  dataKnown_3 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  dataKnown_4 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  dataKnown_5 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  dataKnown_6 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  dataKnown_7 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  loadCompleted_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  loadCompleted_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  loadCompleted_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  loadCompleted_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  loadCompleted_4 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  loadCompleted_5 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  loadCompleted_6 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  loadCompleted_7 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  bypassInitiated_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  bypassInitiated_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  bypassInitiated_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  bypassInitiated_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  bypassInitiated_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  bypassInitiated_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  bypassInitiated_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  bypassInitiated_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  checkBits_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  checkBits_1 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  checkBits_2 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  checkBits_3 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  checkBits_4 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  checkBits_5 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  checkBits_6 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  checkBits_7 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  previousStoreHead = _RAND_82[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  conflictPReg_0_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  conflictPReg_0_1 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  conflictPReg_0_2 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  conflictPReg_0_3 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  conflictPReg_0_4 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  conflictPReg_0_5 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  conflictPReg_0_6 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  conflictPReg_0_7 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  conflictPReg_1_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  conflictPReg_1_1 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  conflictPReg_1_2 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  conflictPReg_1_3 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  conflictPReg_1_4 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  conflictPReg_1_5 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  conflictPReg_1_6 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  conflictPReg_1_7 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  conflictPReg_2_0 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  conflictPReg_2_1 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  conflictPReg_2_2 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  conflictPReg_2_3 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  conflictPReg_2_4 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  conflictPReg_2_5 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  conflictPReg_2_6 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  conflictPReg_2_7 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  conflictPReg_3_0 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  conflictPReg_3_1 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  conflictPReg_3_2 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  conflictPReg_3_3 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  conflictPReg_3_4 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  conflictPReg_3_5 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  conflictPReg_3_6 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  conflictPReg_3_7 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  conflictPReg_4_0 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  conflictPReg_4_1 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  conflictPReg_4_2 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  conflictPReg_4_3 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  conflictPReg_4_4 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  conflictPReg_4_5 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  conflictPReg_4_6 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  conflictPReg_4_7 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  conflictPReg_5_0 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  conflictPReg_5_1 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  conflictPReg_5_2 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  conflictPReg_5_3 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  conflictPReg_5_4 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  conflictPReg_5_5 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  conflictPReg_5_6 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  conflictPReg_5_7 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  conflictPReg_6_0 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  conflictPReg_6_1 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  conflictPReg_6_2 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  conflictPReg_6_3 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  conflictPReg_6_4 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  conflictPReg_6_5 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  conflictPReg_6_6 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  conflictPReg_6_7 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  conflictPReg_7_0 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  conflictPReg_7_1 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  conflictPReg_7_2 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  conflictPReg_7_3 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  conflictPReg_7_4 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  conflictPReg_7_5 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  conflictPReg_7_6 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  conflictPReg_7_7 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_0 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_1 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_2 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_3 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_4 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_5 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_6 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_7 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_0 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_1 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_2 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_3 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_4 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_5 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_6 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_7 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_0 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_1 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_2 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_3 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_4 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_5 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_6 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_7 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_0 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_1 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_2 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_3 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_4 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_5 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_6 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_7 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_0 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_1 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_2 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_3 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_4 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_5 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_6 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_7 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_0 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_1 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_2 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_3 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_4 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_5 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_6 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_7 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_0 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_1 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_2 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_3 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_4 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_5 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_6 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_7 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_0 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_1 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_2 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_3 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_4 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_5 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_6 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_7 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_0 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_1 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_2 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_3 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_4 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_5 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_6 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_7 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  shiftedStoreDataQPreg_0 = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  shiftedStoreDataQPreg_1 = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  shiftedStoreDataQPreg_2 = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  shiftedStoreDataQPreg_3 = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  shiftedStoreDataQPreg_4 = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  shiftedStoreDataQPreg_5 = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  shiftedStoreDataQPreg_6 = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  shiftedStoreDataQPreg_7 = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  addrKnownPReg_0 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  addrKnownPReg_1 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  addrKnownPReg_2 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  addrKnownPReg_3 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  addrKnownPReg_4 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  addrKnownPReg_5 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  addrKnownPReg_6 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  addrKnownPReg_7 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  dataKnownPReg_0 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  dataKnownPReg_1 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  dataKnownPReg_2 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  dataKnownPReg_3 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  dataKnownPReg_4 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  dataKnownPReg_5 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  dataKnownPReg_6 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  dataKnownPReg_7 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  prevPriorityRequest_7 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  prevPriorityRequest_6 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  prevPriorityRequest_5 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  prevPriorityRequest_4 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  prevPriorityRequest_3 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  prevPriorityRequest_2 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  prevPriorityRequest_1 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  prevPriorityRequest_0 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 3'h0;
    end else begin
      head <= _GEN_764[2:0];
    end
    if (reset) begin
      tail <= 3'h0;
    end else begin
      tail <= _GEN_765[2:0];
    end
    if (reset) begin
      offsetQ_0 <= 3'h0;
    end else begin
      if (initBits_0) begin
        if (3'h7 == _T_1156) begin
          offsetQ_0 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1156) begin
            offsetQ_0 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1156) begin
              offsetQ_0 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1156) begin
                offsetQ_0 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1156) begin
                  offsetQ_0 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1156) begin
                    offsetQ_0 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1156) begin
                      offsetQ_0 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_0 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 3'h0;
    end else begin
      if (initBits_1) begin
        if (3'h7 == _T_1174) begin
          offsetQ_1 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1174) begin
            offsetQ_1 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1174) begin
              offsetQ_1 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1174) begin
                offsetQ_1 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1174) begin
                  offsetQ_1 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1174) begin
                    offsetQ_1 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1174) begin
                      offsetQ_1 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_1 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 3'h0;
    end else begin
      if (initBits_2) begin
        if (3'h7 == _T_1192) begin
          offsetQ_2 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1192) begin
            offsetQ_2 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1192) begin
              offsetQ_2 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1192) begin
                offsetQ_2 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1192) begin
                  offsetQ_2 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1192) begin
                    offsetQ_2 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1192) begin
                      offsetQ_2 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_2 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 3'h0;
    end else begin
      if (initBits_3) begin
        if (3'h7 == _T_1210) begin
          offsetQ_3 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1210) begin
            offsetQ_3 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1210) begin
              offsetQ_3 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1210) begin
                offsetQ_3 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1210) begin
                  offsetQ_3 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1210) begin
                    offsetQ_3 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1210) begin
                      offsetQ_3 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_3 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 3'h0;
    end else begin
      if (initBits_4) begin
        if (3'h7 == _T_1228) begin
          offsetQ_4 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1228) begin
            offsetQ_4 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1228) begin
              offsetQ_4 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1228) begin
                offsetQ_4 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1228) begin
                  offsetQ_4 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1228) begin
                    offsetQ_4 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1228) begin
                      offsetQ_4 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_4 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 3'h0;
    end else begin
      if (initBits_5) begin
        if (3'h7 == _T_1246) begin
          offsetQ_5 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1246) begin
            offsetQ_5 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1246) begin
              offsetQ_5 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1246) begin
                offsetQ_5 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1246) begin
                  offsetQ_5 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1246) begin
                    offsetQ_5 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1246) begin
                      offsetQ_5 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_5 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 3'h0;
    end else begin
      if (initBits_6) begin
        if (3'h7 == _T_1264) begin
          offsetQ_6 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1264) begin
            offsetQ_6 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1264) begin
              offsetQ_6 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1264) begin
                offsetQ_6 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1264) begin
                  offsetQ_6 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1264) begin
                    offsetQ_6 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1264) begin
                      offsetQ_6 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_6 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 3'h0;
    end else begin
      if (initBits_7) begin
        if (3'h7 == _T_1282) begin
          offsetQ_7 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1282) begin
            offsetQ_7 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1282) begin
              offsetQ_7 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1282) begin
                offsetQ_7 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1282) begin
                  offsetQ_7 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1282) begin
                    offsetQ_7 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1282) begin
                      offsetQ_7 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_7 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 3'h0;
    end else begin
      if (initBits_0) begin
        if (3'h7 == _T_1156) begin
          portQ_0 <= 3'h0;
        end else begin
          if (3'h6 == _T_1156) begin
            portQ_0 <= 3'h0;
          end else begin
            if (3'h5 == _T_1156) begin
              portQ_0 <= 3'h0;
            end else begin
              if (3'h4 == _T_1156) begin
                portQ_0 <= 3'h0;
              end else begin
                if (3'h3 == _T_1156) begin
                  portQ_0 <= 3'h0;
                end else begin
                  if (3'h2 == _T_1156) begin
                    portQ_0 <= io_bbLoadPorts_2;
                  end else begin
                    if (3'h1 == _T_1156) begin
                      portQ_0 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_0 <= io_bbLoadPorts_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_1 <= 3'h0;
    end else begin
      if (initBits_1) begin
        if (3'h7 == _T_1174) begin
          portQ_1 <= 3'h0;
        end else begin
          if (3'h6 == _T_1174) begin
            portQ_1 <= 3'h0;
          end else begin
            if (3'h5 == _T_1174) begin
              portQ_1 <= 3'h0;
            end else begin
              if (3'h4 == _T_1174) begin
                portQ_1 <= 3'h0;
              end else begin
                if (3'h3 == _T_1174) begin
                  portQ_1 <= 3'h0;
                end else begin
                  if (3'h2 == _T_1174) begin
                    portQ_1 <= io_bbLoadPorts_2;
                  end else begin
                    if (3'h1 == _T_1174) begin
                      portQ_1 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_1 <= io_bbLoadPorts_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_2 <= 3'h0;
    end else begin
      if (initBits_2) begin
        if (3'h7 == _T_1192) begin
          portQ_2 <= 3'h0;
        end else begin
          if (3'h6 == _T_1192) begin
            portQ_2 <= 3'h0;
          end else begin
            if (3'h5 == _T_1192) begin
              portQ_2 <= 3'h0;
            end else begin
              if (3'h4 == _T_1192) begin
                portQ_2 <= 3'h0;
              end else begin
                if (3'h3 == _T_1192) begin
                  portQ_2 <= 3'h0;
                end else begin
                  if (3'h2 == _T_1192) begin
                    portQ_2 <= io_bbLoadPorts_2;
                  end else begin
                    if (3'h1 == _T_1192) begin
                      portQ_2 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_2 <= io_bbLoadPorts_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_3 <= 3'h0;
    end else begin
      if (initBits_3) begin
        if (3'h7 == _T_1210) begin
          portQ_3 <= 3'h0;
        end else begin
          if (3'h6 == _T_1210) begin
            portQ_3 <= 3'h0;
          end else begin
            if (3'h5 == _T_1210) begin
              portQ_3 <= 3'h0;
            end else begin
              if (3'h4 == _T_1210) begin
                portQ_3 <= 3'h0;
              end else begin
                if (3'h3 == _T_1210) begin
                  portQ_3 <= 3'h0;
                end else begin
                  if (3'h2 == _T_1210) begin
                    portQ_3 <= io_bbLoadPorts_2;
                  end else begin
                    if (3'h1 == _T_1210) begin
                      portQ_3 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_3 <= io_bbLoadPorts_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_4 <= 3'h0;
    end else begin
      if (initBits_4) begin
        if (3'h7 == _T_1228) begin
          portQ_4 <= 3'h0;
        end else begin
          if (3'h6 == _T_1228) begin
            portQ_4 <= 3'h0;
          end else begin
            if (3'h5 == _T_1228) begin
              portQ_4 <= 3'h0;
            end else begin
              if (3'h4 == _T_1228) begin
                portQ_4 <= 3'h0;
              end else begin
                if (3'h3 == _T_1228) begin
                  portQ_4 <= 3'h0;
                end else begin
                  if (3'h2 == _T_1228) begin
                    portQ_4 <= io_bbLoadPorts_2;
                  end else begin
                    if (3'h1 == _T_1228) begin
                      portQ_4 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_4 <= io_bbLoadPorts_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_5 <= 3'h0;
    end else begin
      if (initBits_5) begin
        if (3'h7 == _T_1246) begin
          portQ_5 <= 3'h0;
        end else begin
          if (3'h6 == _T_1246) begin
            portQ_5 <= 3'h0;
          end else begin
            if (3'h5 == _T_1246) begin
              portQ_5 <= 3'h0;
            end else begin
              if (3'h4 == _T_1246) begin
                portQ_5 <= 3'h0;
              end else begin
                if (3'h3 == _T_1246) begin
                  portQ_5 <= 3'h0;
                end else begin
                  if (3'h2 == _T_1246) begin
                    portQ_5 <= io_bbLoadPorts_2;
                  end else begin
                    if (3'h1 == _T_1246) begin
                      portQ_5 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_5 <= io_bbLoadPorts_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_6 <= 3'h0;
    end else begin
      if (initBits_6) begin
        if (3'h7 == _T_1264) begin
          portQ_6 <= 3'h0;
        end else begin
          if (3'h6 == _T_1264) begin
            portQ_6 <= 3'h0;
          end else begin
            if (3'h5 == _T_1264) begin
              portQ_6 <= 3'h0;
            end else begin
              if (3'h4 == _T_1264) begin
                portQ_6 <= 3'h0;
              end else begin
                if (3'h3 == _T_1264) begin
                  portQ_6 <= 3'h0;
                end else begin
                  if (3'h2 == _T_1264) begin
                    portQ_6 <= io_bbLoadPorts_2;
                  end else begin
                    if (3'h1 == _T_1264) begin
                      portQ_6 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_6 <= io_bbLoadPorts_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_7 <= 3'h0;
    end else begin
      if (initBits_7) begin
        if (3'h7 == _T_1282) begin
          portQ_7 <= 3'h0;
        end else begin
          if (3'h6 == _T_1282) begin
            portQ_7 <= 3'h0;
          end else begin
            if (3'h5 == _T_1282) begin
              portQ_7 <= 3'h0;
            end else begin
              if (3'h4 == _T_1282) begin
                portQ_7 <= 3'h0;
              end else begin
                if (3'h3 == _T_1282) begin
                  portQ_7 <= 3'h0;
                end else begin
                  if (3'h2 == _T_1282) begin
                    portQ_7 <= io_bbLoadPorts_2;
                  end else begin
                    if (3'h1 == _T_1282) begin
                      portQ_7 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_7 <= io_bbLoadPorts_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_31522) begin
          if (3'h4 == _T_31539) begin
            addrQ_0 <= io_addrFromLoadPorts_4;
          end else begin
            if (3'h3 == _T_31539) begin
              addrQ_0 <= io_addrFromLoadPorts_3;
            end else begin
              if (3'h2 == _T_31539) begin
                addrQ_0 <= io_addrFromLoadPorts_2;
              end else begin
                if (3'h1 == _T_31539) begin
                  addrQ_0 <= io_addrFromLoadPorts_1;
                end else begin
                  addrQ_0 <= io_addrFromLoadPorts_0;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_31564) begin
          if (3'h4 == _T_31581) begin
            addrQ_1 <= io_addrFromLoadPorts_4;
          end else begin
            if (3'h3 == _T_31581) begin
              addrQ_1 <= io_addrFromLoadPorts_3;
            end else begin
              if (3'h2 == _T_31581) begin
                addrQ_1 <= io_addrFromLoadPorts_2;
              end else begin
                if (3'h1 == _T_31581) begin
                  addrQ_1 <= io_addrFromLoadPorts_1;
                end else begin
                  addrQ_1 <= io_addrFromLoadPorts_0;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_31606) begin
          if (3'h4 == _T_31623) begin
            addrQ_2 <= io_addrFromLoadPorts_4;
          end else begin
            if (3'h3 == _T_31623) begin
              addrQ_2 <= io_addrFromLoadPorts_3;
            end else begin
              if (3'h2 == _T_31623) begin
                addrQ_2 <= io_addrFromLoadPorts_2;
              end else begin
                if (3'h1 == _T_31623) begin
                  addrQ_2 <= io_addrFromLoadPorts_1;
                end else begin
                  addrQ_2 <= io_addrFromLoadPorts_0;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_31648) begin
          if (3'h4 == _T_31665) begin
            addrQ_3 <= io_addrFromLoadPorts_4;
          end else begin
            if (3'h3 == _T_31665) begin
              addrQ_3 <= io_addrFromLoadPorts_3;
            end else begin
              if (3'h2 == _T_31665) begin
                addrQ_3 <= io_addrFromLoadPorts_2;
              end else begin
                if (3'h1 == _T_31665) begin
                  addrQ_3 <= io_addrFromLoadPorts_1;
                end else begin
                  addrQ_3 <= io_addrFromLoadPorts_0;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_31690) begin
          if (3'h4 == _T_31707) begin
            addrQ_4 <= io_addrFromLoadPorts_4;
          end else begin
            if (3'h3 == _T_31707) begin
              addrQ_4 <= io_addrFromLoadPorts_3;
            end else begin
              if (3'h2 == _T_31707) begin
                addrQ_4 <= io_addrFromLoadPorts_2;
              end else begin
                if (3'h1 == _T_31707) begin
                  addrQ_4 <= io_addrFromLoadPorts_1;
                end else begin
                  addrQ_4 <= io_addrFromLoadPorts_0;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_31732) begin
          if (3'h4 == _T_31749) begin
            addrQ_5 <= io_addrFromLoadPorts_4;
          end else begin
            if (3'h3 == _T_31749) begin
              addrQ_5 <= io_addrFromLoadPorts_3;
            end else begin
              if (3'h2 == _T_31749) begin
                addrQ_5 <= io_addrFromLoadPorts_2;
              end else begin
                if (3'h1 == _T_31749) begin
                  addrQ_5 <= io_addrFromLoadPorts_1;
                end else begin
                  addrQ_5 <= io_addrFromLoadPorts_0;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_31774) begin
          if (3'h4 == _T_31791) begin
            addrQ_6 <= io_addrFromLoadPorts_4;
          end else begin
            if (3'h3 == _T_31791) begin
              addrQ_6 <= io_addrFromLoadPorts_3;
            end else begin
              if (3'h2 == _T_31791) begin
                addrQ_6 <= io_addrFromLoadPorts_2;
              end else begin
                if (3'h1 == _T_31791) begin
                  addrQ_6 <= io_addrFromLoadPorts_1;
                end else begin
                  addrQ_6 <= io_addrFromLoadPorts_0;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_31816) begin
          if (3'h4 == _T_31833) begin
            addrQ_7 <= io_addrFromLoadPorts_4;
          end else begin
            if (3'h3 == _T_31833) begin
              addrQ_7 <= io_addrFromLoadPorts_3;
            end else begin
              if (3'h2 == _T_31833) begin
                addrQ_7 <= io_addrFromLoadPorts_2;
              end else begin
                if (3'h1 == _T_31833) begin
                  addrQ_7 <= io_addrFromLoadPorts_1;
                end else begin
                  addrQ_7 <= io_addrFromLoadPorts_0;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (bypassRequest_0) begin
        if (_T_23570) begin
          if (3'h7 == _T_23561) begin
            dataQ_0 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23561) begin
              dataQ_0 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23561) begin
                dataQ_0 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23561) begin
                  dataQ_0 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23561) begin
                    dataQ_0 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23561) begin
                      dataQ_0 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23561) begin
                        dataQ_0 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_0 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_0 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_0) begin
          dataQ_0 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (bypassRequest_1) begin
        if (_T_23650) begin
          if (3'h7 == _T_23641) begin
            dataQ_1 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23641) begin
              dataQ_1 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23641) begin
                dataQ_1 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23641) begin
                  dataQ_1 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23641) begin
                    dataQ_1 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23641) begin
                      dataQ_1 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23641) begin
                        dataQ_1 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_1 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_1 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_1) begin
          dataQ_1 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (bypassRequest_2) begin
        if (_T_23730) begin
          if (3'h7 == _T_23721) begin
            dataQ_2 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23721) begin
              dataQ_2 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23721) begin
                dataQ_2 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23721) begin
                  dataQ_2 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23721) begin
                    dataQ_2 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23721) begin
                      dataQ_2 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23721) begin
                        dataQ_2 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_2 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_2 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_2) begin
          dataQ_2 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (bypassRequest_3) begin
        if (_T_23810) begin
          if (3'h7 == _T_23801) begin
            dataQ_3 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23801) begin
              dataQ_3 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23801) begin
                dataQ_3 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23801) begin
                  dataQ_3 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23801) begin
                    dataQ_3 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23801) begin
                      dataQ_3 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23801) begin
                        dataQ_3 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_3 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_3 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_3) begin
          dataQ_3 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (bypassRequest_4) begin
        if (_T_23890) begin
          if (3'h7 == _T_23881) begin
            dataQ_4 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23881) begin
              dataQ_4 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23881) begin
                dataQ_4 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23881) begin
                  dataQ_4 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23881) begin
                    dataQ_4 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23881) begin
                      dataQ_4 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23881) begin
                        dataQ_4 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_4 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_4 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_4) begin
          dataQ_4 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (bypassRequest_5) begin
        if (_T_23970) begin
          if (3'h7 == _T_23961) begin
            dataQ_5 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23961) begin
              dataQ_5 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23961) begin
                dataQ_5 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23961) begin
                  dataQ_5 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23961) begin
                    dataQ_5 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23961) begin
                      dataQ_5 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23961) begin
                        dataQ_5 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_5 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_5 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_5) begin
          dataQ_5 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (bypassRequest_6) begin
        if (_T_24050) begin
          if (3'h7 == _T_24041) begin
            dataQ_6 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_24041) begin
              dataQ_6 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_24041) begin
                dataQ_6 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_24041) begin
                  dataQ_6 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_24041) begin
                    dataQ_6 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_24041) begin
                      dataQ_6 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_24041) begin
                        dataQ_6 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_6 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_6 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_6) begin
          dataQ_6 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (bypassRequest_7) begin
        if (_T_24130) begin
          if (3'h7 == _T_24121) begin
            dataQ_7 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_24121) begin
              dataQ_7 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_24121) begin
                dataQ_7 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_24121) begin
                  dataQ_7 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_24121) begin
                    dataQ_7 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_24121) begin
                      dataQ_7 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_24121) begin
                        dataQ_7 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_7 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_7 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_7) begin
          dataQ_7 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_31522) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_31564) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_31606) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_31648) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_31690) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_31732) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_31774) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_31816) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_25249) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_25252) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_25255) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_25258) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_25261) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_25264) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_25267) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_25270) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        loadCompleted_0 <= 1'h0;
      end else begin
        if (loadCompleting_0) begin
          loadCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        loadCompleted_1 <= 1'h0;
      end else begin
        if (loadCompleting_1) begin
          loadCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        loadCompleted_2 <= 1'h0;
      end else begin
        if (loadCompleting_2) begin
          loadCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        loadCompleted_3 <= 1'h0;
      end else begin
        if (loadCompleting_3) begin
          loadCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        loadCompleted_4 <= 1'h0;
      end else begin
        if (loadCompleting_4) begin
          loadCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        loadCompleted_5 <= 1'h0;
      end else begin
        if (loadCompleting_5) begin
          loadCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        loadCompleted_6 <= 1'h0;
      end else begin
        if (loadCompleting_6) begin
          loadCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        loadCompleted_7 <= 1'h0;
      end else begin
        if (loadCompleting_7) begin
          loadCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1126;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1127;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1128;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1129;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1130;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1131;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1132;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1133;
    end
    if (reset) begin
      bypassInitiated_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        bypassInitiated_0 <= 1'h0;
      end else begin
        if (bypassRequest_0) begin
          bypassInitiated_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        bypassInitiated_1 <= 1'h0;
      end else begin
        if (bypassRequest_1) begin
          bypassInitiated_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        bypassInitiated_2 <= 1'h0;
      end else begin
        if (bypassRequest_2) begin
          bypassInitiated_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        bypassInitiated_3 <= 1'h0;
      end else begin
        if (bypassRequest_3) begin
          bypassInitiated_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        bypassInitiated_4 <= 1'h0;
      end else begin
        if (bypassRequest_4) begin
          bypassInitiated_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        bypassInitiated_5 <= 1'h0;
      end else begin
        if (bypassRequest_5) begin
          bypassInitiated_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        bypassInitiated_6 <= 1'h0;
      end else begin
        if (bypassRequest_6) begin
          bypassInitiated_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        bypassInitiated_7 <= 1'h0;
      end else begin
        if (bypassRequest_7) begin
          bypassInitiated_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_1309;
      end else begin
        if (io_storeEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_1313) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_1321) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_1339;
      end else begin
        if (io_storeEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_1343) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_1351) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_1369;
      end else begin
        if (io_storeEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_1373) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_1381) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_1399;
      end else begin
        if (io_storeEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_1403) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_1411) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_1429;
      end else begin
        if (io_storeEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_1433) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_1441) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_1459;
      end else begin
        if (io_storeEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_1463) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_1471) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_1489;
      end else begin
        if (io_storeEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_1493) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_1501) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_1519;
      end else begin
        if (io_storeEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_1523) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_1531) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    previousStoreHead <= io_storeHead;
    conflictPReg_0_0 <= _T_6218[0];
    conflictPReg_0_1 <= _T_6218[1];
    conflictPReg_0_2 <= _T_6218[2];
    conflictPReg_0_3 <= _T_6218[3];
    conflictPReg_0_4 <= _T_6218[4];
    conflictPReg_0_5 <= _T_6218[5];
    conflictPReg_0_6 <= _T_6218[6];
    conflictPReg_0_7 <= _T_6218[7];
    conflictPReg_1_0 <= _T_6532[0];
    conflictPReg_1_1 <= _T_6532[1];
    conflictPReg_1_2 <= _T_6532[2];
    conflictPReg_1_3 <= _T_6532[3];
    conflictPReg_1_4 <= _T_6532[4];
    conflictPReg_1_5 <= _T_6532[5];
    conflictPReg_1_6 <= _T_6532[6];
    conflictPReg_1_7 <= _T_6532[7];
    conflictPReg_2_0 <= _T_6846[0];
    conflictPReg_2_1 <= _T_6846[1];
    conflictPReg_2_2 <= _T_6846[2];
    conflictPReg_2_3 <= _T_6846[3];
    conflictPReg_2_4 <= _T_6846[4];
    conflictPReg_2_5 <= _T_6846[5];
    conflictPReg_2_6 <= _T_6846[6];
    conflictPReg_2_7 <= _T_6846[7];
    conflictPReg_3_0 <= _T_7160[0];
    conflictPReg_3_1 <= _T_7160[1];
    conflictPReg_3_2 <= _T_7160[2];
    conflictPReg_3_3 <= _T_7160[3];
    conflictPReg_3_4 <= _T_7160[4];
    conflictPReg_3_5 <= _T_7160[5];
    conflictPReg_3_6 <= _T_7160[6];
    conflictPReg_3_7 <= _T_7160[7];
    conflictPReg_4_0 <= _T_7474[0];
    conflictPReg_4_1 <= _T_7474[1];
    conflictPReg_4_2 <= _T_7474[2];
    conflictPReg_4_3 <= _T_7474[3];
    conflictPReg_4_4 <= _T_7474[4];
    conflictPReg_4_5 <= _T_7474[5];
    conflictPReg_4_6 <= _T_7474[6];
    conflictPReg_4_7 <= _T_7474[7];
    conflictPReg_5_0 <= _T_7788[0];
    conflictPReg_5_1 <= _T_7788[1];
    conflictPReg_5_2 <= _T_7788[2];
    conflictPReg_5_3 <= _T_7788[3];
    conflictPReg_5_4 <= _T_7788[4];
    conflictPReg_5_5 <= _T_7788[5];
    conflictPReg_5_6 <= _T_7788[6];
    conflictPReg_5_7 <= _T_7788[7];
    conflictPReg_6_0 <= _T_8102[0];
    conflictPReg_6_1 <= _T_8102[1];
    conflictPReg_6_2 <= _T_8102[2];
    conflictPReg_6_3 <= _T_8102[3];
    conflictPReg_6_4 <= _T_8102[4];
    conflictPReg_6_5 <= _T_8102[5];
    conflictPReg_6_6 <= _T_8102[6];
    conflictPReg_6_7 <= _T_8102[7];
    conflictPReg_7_0 <= _T_8416[0];
    conflictPReg_7_1 <= _T_8416[1];
    conflictPReg_7_2 <= _T_8416[2];
    conflictPReg_7_3 <= _T_8416[3];
    conflictPReg_7_4 <= _T_8416[4];
    conflictPReg_7_5 <= _T_8416[5];
    conflictPReg_7_6 <= _T_8416[6];
    conflictPReg_7_7 <= _T_8416[7];
    storeAddrNotKnownFlagsPReg_0_0 <= _T_14598[0];
    storeAddrNotKnownFlagsPReg_0_1 <= _T_14598[1];
    storeAddrNotKnownFlagsPReg_0_2 <= _T_14598[2];
    storeAddrNotKnownFlagsPReg_0_3 <= _T_14598[3];
    storeAddrNotKnownFlagsPReg_0_4 <= _T_14598[4];
    storeAddrNotKnownFlagsPReg_0_5 <= _T_14598[5];
    storeAddrNotKnownFlagsPReg_0_6 <= _T_14598[6];
    storeAddrNotKnownFlagsPReg_0_7 <= _T_14598[7];
    storeAddrNotKnownFlagsPReg_1_0 <= _T_14912[0];
    storeAddrNotKnownFlagsPReg_1_1 <= _T_14912[1];
    storeAddrNotKnownFlagsPReg_1_2 <= _T_14912[2];
    storeAddrNotKnownFlagsPReg_1_3 <= _T_14912[3];
    storeAddrNotKnownFlagsPReg_1_4 <= _T_14912[4];
    storeAddrNotKnownFlagsPReg_1_5 <= _T_14912[5];
    storeAddrNotKnownFlagsPReg_1_6 <= _T_14912[6];
    storeAddrNotKnownFlagsPReg_1_7 <= _T_14912[7];
    storeAddrNotKnownFlagsPReg_2_0 <= _T_15226[0];
    storeAddrNotKnownFlagsPReg_2_1 <= _T_15226[1];
    storeAddrNotKnownFlagsPReg_2_2 <= _T_15226[2];
    storeAddrNotKnownFlagsPReg_2_3 <= _T_15226[3];
    storeAddrNotKnownFlagsPReg_2_4 <= _T_15226[4];
    storeAddrNotKnownFlagsPReg_2_5 <= _T_15226[5];
    storeAddrNotKnownFlagsPReg_2_6 <= _T_15226[6];
    storeAddrNotKnownFlagsPReg_2_7 <= _T_15226[7];
    storeAddrNotKnownFlagsPReg_3_0 <= _T_15540[0];
    storeAddrNotKnownFlagsPReg_3_1 <= _T_15540[1];
    storeAddrNotKnownFlagsPReg_3_2 <= _T_15540[2];
    storeAddrNotKnownFlagsPReg_3_3 <= _T_15540[3];
    storeAddrNotKnownFlagsPReg_3_4 <= _T_15540[4];
    storeAddrNotKnownFlagsPReg_3_5 <= _T_15540[5];
    storeAddrNotKnownFlagsPReg_3_6 <= _T_15540[6];
    storeAddrNotKnownFlagsPReg_3_7 <= _T_15540[7];
    storeAddrNotKnownFlagsPReg_4_0 <= _T_15854[0];
    storeAddrNotKnownFlagsPReg_4_1 <= _T_15854[1];
    storeAddrNotKnownFlagsPReg_4_2 <= _T_15854[2];
    storeAddrNotKnownFlagsPReg_4_3 <= _T_15854[3];
    storeAddrNotKnownFlagsPReg_4_4 <= _T_15854[4];
    storeAddrNotKnownFlagsPReg_4_5 <= _T_15854[5];
    storeAddrNotKnownFlagsPReg_4_6 <= _T_15854[6];
    storeAddrNotKnownFlagsPReg_4_7 <= _T_15854[7];
    storeAddrNotKnownFlagsPReg_5_0 <= _T_16168[0];
    storeAddrNotKnownFlagsPReg_5_1 <= _T_16168[1];
    storeAddrNotKnownFlagsPReg_5_2 <= _T_16168[2];
    storeAddrNotKnownFlagsPReg_5_3 <= _T_16168[3];
    storeAddrNotKnownFlagsPReg_5_4 <= _T_16168[4];
    storeAddrNotKnownFlagsPReg_5_5 <= _T_16168[5];
    storeAddrNotKnownFlagsPReg_5_6 <= _T_16168[6];
    storeAddrNotKnownFlagsPReg_5_7 <= _T_16168[7];
    storeAddrNotKnownFlagsPReg_6_0 <= _T_16482[0];
    storeAddrNotKnownFlagsPReg_6_1 <= _T_16482[1];
    storeAddrNotKnownFlagsPReg_6_2 <= _T_16482[2];
    storeAddrNotKnownFlagsPReg_6_3 <= _T_16482[3];
    storeAddrNotKnownFlagsPReg_6_4 <= _T_16482[4];
    storeAddrNotKnownFlagsPReg_6_5 <= _T_16482[5];
    storeAddrNotKnownFlagsPReg_6_6 <= _T_16482[6];
    storeAddrNotKnownFlagsPReg_6_7 <= _T_16482[7];
    storeAddrNotKnownFlagsPReg_7_0 <= _T_16796[0];
    storeAddrNotKnownFlagsPReg_7_1 <= _T_16796[1];
    storeAddrNotKnownFlagsPReg_7_2 <= _T_16796[2];
    storeAddrNotKnownFlagsPReg_7_3 <= _T_16796[3];
    storeAddrNotKnownFlagsPReg_7_4 <= _T_16796[4];
    storeAddrNotKnownFlagsPReg_7_5 <= _T_16796[5];
    storeAddrNotKnownFlagsPReg_7_6 <= _T_16796[6];
    storeAddrNotKnownFlagsPReg_7_7 <= _T_16796[7];
    shiftedStoreDataKnownPReg_0 <= _T_2708[0];
    shiftedStoreDataKnownPReg_1 <= _T_2708[1];
    shiftedStoreDataKnownPReg_2 <= _T_2708[2];
    shiftedStoreDataKnownPReg_3 <= _T_2708[3];
    shiftedStoreDataKnownPReg_4 <= _T_2708[4];
    shiftedStoreDataKnownPReg_5 <= _T_2708[5];
    shiftedStoreDataKnownPReg_6 <= _T_2708[6];
    shiftedStoreDataKnownPReg_7 <= _T_2708[7];
    shiftedStoreDataQPreg_0 <= _T_2395[31:0];
    shiftedStoreDataQPreg_1 <= _T_2395[63:32];
    shiftedStoreDataQPreg_2 <= _T_2395[95:64];
    shiftedStoreDataQPreg_3 <= _T_2395[127:96];
    shiftedStoreDataQPreg_4 <= _T_2395[159:128];
    shiftedStoreDataQPreg_5 <= _T_2395[191:160];
    shiftedStoreDataQPreg_6 <= _T_2395[223:192];
    shiftedStoreDataQPreg_7 <= _T_2395[255:224];
    addrKnownPReg_0 <= addrKnown_0;
    addrKnownPReg_1 <= addrKnown_1;
    addrKnownPReg_2 <= addrKnown_2;
    addrKnownPReg_3 <= addrKnown_3;
    addrKnownPReg_4 <= addrKnown_4;
    addrKnownPReg_5 <= addrKnown_5;
    addrKnownPReg_6 <= addrKnown_6;
    addrKnownPReg_7 <= addrKnown_7;
    dataKnownPReg_0 <= dataKnown_0;
    dataKnownPReg_1 <= dataKnown_1;
    dataKnownPReg_2 <= dataKnown_2;
    dataKnownPReg_3 <= dataKnown_3;
    dataKnownPReg_4 <= dataKnown_4;
    dataKnownPReg_5 <= dataKnown_5;
    dataKnownPReg_6 <= dataKnown_6;
    dataKnownPReg_7 <= dataKnown_7;
    if (reset) begin
      prevPriorityRequest_7 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_7 <= priorityLoadRequest_7;
      end else begin
        prevPriorityRequest_7 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_6 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_6 <= priorityLoadRequest_6;
      end else begin
        prevPriorityRequest_6 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_5 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_5 <= priorityLoadRequest_5;
      end else begin
        prevPriorityRequest_5 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_4 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_4 <= priorityLoadRequest_4;
      end else begin
        prevPriorityRequest_4 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_3 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_3 <= priorityLoadRequest_3;
      end else begin
        prevPriorityRequest_3 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_2 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_2 <= priorityLoadRequest_2;
      end else begin
        prevPriorityRequest_2 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_1 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_1 <= priorityLoadRequest_1;
      end else begin
        prevPriorityRequest_1 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_0 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_0 <= priorityLoadRequest_0;
      end else begin
        prevPriorityRequest_0 <= 1'h0;
      end
    end
  end
endmodule
module GROUP_ALLOCATOR_LSQ_dist( // @[:@13723.2]
  output [2:0] io_bbLoadOffsets_0, // @[:@13726.4]
  output [2:0] io_bbLoadOffsets_1, // @[:@13726.4]
  output [2:0] io_bbLoadOffsets_2, // @[:@13726.4]
  output [2:0] io_bbLoadOffsets_3, // @[:@13726.4]
  output [2:0] io_bbLoadOffsets_4, // @[:@13726.4]
  output [2:0] io_bbLoadOffsets_5, // @[:@13726.4]
  output [2:0] io_bbLoadOffsets_6, // @[:@13726.4]
  output [2:0] io_bbLoadOffsets_7, // @[:@13726.4]
  output [2:0] io_bbLoadPorts_0, // @[:@13726.4]
  output [2:0] io_bbLoadPorts_1, // @[:@13726.4]
  output [2:0] io_bbLoadPorts_2, // @[:@13726.4]
  output [2:0] io_bbNumLoads, // @[:@13726.4]
  input  [2:0] io_loadTail, // @[:@13726.4]
  input  [2:0] io_loadHead, // @[:@13726.4]
  input        io_loadEmpty, // @[:@13726.4]
  output [2:0] io_bbStoreOffsets_0, // @[:@13726.4]
  output [2:0] io_bbStoreOffsets_1, // @[:@13726.4]
  output [2:0] io_bbStoreOffsets_2, // @[:@13726.4]
  output [2:0] io_bbStoreOffsets_3, // @[:@13726.4]
  output [2:0] io_bbStoreOffsets_4, // @[:@13726.4]
  output [2:0] io_bbStoreOffsets_5, // @[:@13726.4]
  output [2:0] io_bbStoreOffsets_6, // @[:@13726.4]
  output [2:0] io_bbStoreOffsets_7, // @[:@13726.4]
  output       io_bbNumStores, // @[:@13726.4]
  input  [2:0] io_storeTail, // @[:@13726.4]
  input  [2:0] io_storeHead, // @[:@13726.4]
  input        io_storeEmpty, // @[:@13726.4]
  output       io_bbStart, // @[:@13726.4]
  input        io_bbStartSignals_0, // @[:@13726.4]
  input        io_bbStartSignals_1, // @[:@13726.4]
  output       io_readyToPrevious_0, // @[:@13726.4]
  output       io_readyToPrevious_1, // @[:@13726.4]
  output       io_loadPortsEnable_0, // @[:@13726.4]
  output       io_loadPortsEnable_1, // @[:@13726.4]
  output       io_loadPortsEnable_2, // @[:@13726.4]
  output       io_loadPortsEnable_3, // @[:@13726.4]
  output       io_loadPortsEnable_4, // @[:@13726.4]
  output       io_storePortsEnable_0 // @[:@13726.4]
);
  wire  _T_188; // @[GroupAllocator.scala 42:25:@13729.4]
  wire  _T_189; // @[GroupAllocator.scala 42:16:@13730.4]
  wire [3:0] _GEN_36; // @[GroupAllocator.scala 43:36:@13732.6]
  wire [4:0] _T_191; // @[GroupAllocator.scala 43:36:@13732.6]
  wire [4:0] _T_192; // @[GroupAllocator.scala 43:36:@13733.6]
  wire [3:0] _T_193; // @[GroupAllocator.scala 43:36:@13734.6]
  wire [3:0] _GEN_37; // @[GroupAllocator.scala 43:43:@13735.6]
  wire [4:0] _T_194; // @[GroupAllocator.scala 43:43:@13735.6]
  wire [3:0] _T_195; // @[GroupAllocator.scala 43:43:@13736.6]
  wire [3:0] _T_196; // @[GroupAllocator.scala 45:22:@13740.6]
  wire [3:0] _T_197; // @[GroupAllocator.scala 45:22:@13741.6]
  wire [2:0] _T_198; // @[GroupAllocator.scala 45:22:@13742.6]
  wire [3:0] emptyLoadSlots; // @[GroupAllocator.scala 42:34:@13731.4]
  wire  _T_200; // @[GroupAllocator.scala 42:25:@13746.4]
  wire  _T_201; // @[GroupAllocator.scala 42:16:@13747.4]
  wire [3:0] _GEN_38; // @[GroupAllocator.scala 43:36:@13749.6]
  wire [4:0] _T_203; // @[GroupAllocator.scala 43:36:@13749.6]
  wire [4:0] _T_204; // @[GroupAllocator.scala 43:36:@13750.6]
  wire [3:0] _T_205; // @[GroupAllocator.scala 43:36:@13751.6]
  wire [3:0] _GEN_39; // @[GroupAllocator.scala 43:43:@13752.6]
  wire [4:0] _T_206; // @[GroupAllocator.scala 43:43:@13752.6]
  wire [3:0] _T_207; // @[GroupAllocator.scala 43:43:@13753.6]
  wire [3:0] _T_208; // @[GroupAllocator.scala 45:22:@13757.6]
  wire [3:0] _T_209; // @[GroupAllocator.scala 45:22:@13758.6]
  wire [2:0] _T_210; // @[GroupAllocator.scala 45:22:@13759.6]
  wire [3:0] emptyStoreSlots; // @[GroupAllocator.scala 42:34:@13748.4]
  wire  _T_217; // @[GroupAllocator.scala 54:19:@13765.4]
  wire  _T_219; // @[GroupAllocator.scala 54:50:@13766.4]
  wire  possibleAllocations_0; // @[GroupAllocator.scala 56:106:@13773.4]
  wire  possibleAllocations_1; // @[GroupAllocator.scala 56:106:@13774.4]
  wire  allocatedBBIdx; // @[Mux.scala 31:69:@13778.4]
  wire  _T_244; // @[GroupAllocator.scala 69:43:@13782.4]
  wire [1:0] _T_357; // @[Mux.scala 46:16:@13872.6]
  wire [1:0] _T_359; // @[Mux.scala 46:16:@13874.6]
  wire  _T_368; // @[Mux.scala 46:16:@13879.6]
  wire [2:0] _T_438_0; // @[Mux.scala 46:16:@13909.6]
  wire [2:0] _T_438_1; // @[Mux.scala 46:16:@13909.6]
  wire [2:0] _T_459_0; // @[Mux.scala 46:16:@13911.6]
  wire [2:0] _T_459_1; // @[Mux.scala 46:16:@13911.6]
  wire [2:0] _T_459_2; // @[Mux.scala 46:16:@13911.6]
  wire [4:0] _T_614; // @[GroupAllocator.scala 110:34:@13968.6]
  wire [3:0] _T_615; // @[GroupAllocator.scala 110:34:@13969.6]
  wire [4:0] _T_617; // @[GroupAllocator.scala 110:55:@13970.6]
  wire [4:0] _T_618; // @[GroupAllocator.scala 110:55:@13971.6]
  wire [3:0] _T_619; // @[GroupAllocator.scala 110:55:@13972.6]
  wire [4:0] _T_621; // @[util.scala 10:8:@13973.6]
  wire [4:0] _GEN_0; // @[util.scala 10:14:@13974.6]
  wire [3:0] _T_622; // @[util.scala 10:14:@13974.6]
  wire [2:0] _T_752; // @[GroupAllocator.scala 110:90:@14056.6 GroupAllocator.scala 110:90:@14057.6]
  wire [2:0] _T_866_0; // @[Mux.scala 46:16:@14131.6]
  wire [2:0] _T_887_0; // @[Mux.scala 46:16:@14133.6]
  wire [4:0] _T_932; // @[GroupAllocator.scala 115:33:@14151.6]
  wire [3:0] _T_933; // @[GroupAllocator.scala 115:33:@14152.6]
  wire [4:0] _T_935; // @[GroupAllocator.scala 115:54:@14153.6]
  wire [4:0] _T_936; // @[GroupAllocator.scala 115:54:@14154.6]
  wire [3:0] _T_937; // @[GroupAllocator.scala 115:54:@14155.6]
  wire [4:0] _T_939; // @[util.scala 10:8:@14156.6]
  wire [4:0] _GEN_1; // @[util.scala 10:14:@14157.6]
  wire [3:0] _T_940; // @[util.scala 10:14:@14157.6]
  wire [4:0] _T_1066; // @[util.scala 10:8:@14237.6]
  wire [4:0] _GEN_2; // @[util.scala 10:14:@14238.6]
  wire [3:0] _T_1067; // @[util.scala 10:14:@14238.6]
  wire [2:0] _T_1070; // @[GroupAllocator.scala 115:89:@14239.6 GroupAllocator.scala 115:89:@14240.6]
  wire [2:0] _T_1184_0; // @[Mux.scala 46:16:@14314.6]
  wire [2:0] _T_1084; // @[GroupAllocator.scala 115:89:@14248.6 GroupAllocator.scala 115:89:@14249.6]
  wire [2:0] _T_1184_1; // @[Mux.scala 46:16:@14314.6]
  wire [2:0] _T_1205_0; // @[Mux.scala 46:16:@14316.6]
  wire [2:0] _T_1205_1; // @[Mux.scala 46:16:@14316.6]
  assign _T_188 = io_loadHead < io_loadTail; // @[GroupAllocator.scala 42:25:@13729.4]
  assign _T_189 = io_loadEmpty | _T_188; // @[GroupAllocator.scala 42:16:@13730.4]
  assign _GEN_36 = {{1'd0}, io_loadTail}; // @[GroupAllocator.scala 43:36:@13732.6]
  assign _T_191 = 4'h8 - _GEN_36; // @[GroupAllocator.scala 43:36:@13732.6]
  assign _T_192 = $unsigned(_T_191); // @[GroupAllocator.scala 43:36:@13733.6]
  assign _T_193 = _T_192[3:0]; // @[GroupAllocator.scala 43:36:@13734.6]
  assign _GEN_37 = {{1'd0}, io_loadHead}; // @[GroupAllocator.scala 43:43:@13735.6]
  assign _T_194 = _T_193 + _GEN_37; // @[GroupAllocator.scala 43:43:@13735.6]
  assign _T_195 = _T_193 + _GEN_37; // @[GroupAllocator.scala 43:43:@13736.6]
  assign _T_196 = io_loadHead - io_loadTail; // @[GroupAllocator.scala 45:22:@13740.6]
  assign _T_197 = $unsigned(_T_196); // @[GroupAllocator.scala 45:22:@13741.6]
  assign _T_198 = _T_197[2:0]; // @[GroupAllocator.scala 45:22:@13742.6]
  assign emptyLoadSlots = _T_189 ? _T_195 : {{1'd0}, _T_198}; // @[GroupAllocator.scala 42:34:@13731.4]
  assign _T_200 = io_storeHead < io_storeTail; // @[GroupAllocator.scala 42:25:@13746.4]
  assign _T_201 = io_storeEmpty | _T_200; // @[GroupAllocator.scala 42:16:@13747.4]
  assign _GEN_38 = {{1'd0}, io_storeTail}; // @[GroupAllocator.scala 43:36:@13749.6]
  assign _T_203 = 4'h8 - _GEN_38; // @[GroupAllocator.scala 43:36:@13749.6]
  assign _T_204 = $unsigned(_T_203); // @[GroupAllocator.scala 43:36:@13750.6]
  assign _T_205 = _T_204[3:0]; // @[GroupAllocator.scala 43:36:@13751.6]
  assign _GEN_39 = {{1'd0}, io_storeHead}; // @[GroupAllocator.scala 43:43:@13752.6]
  assign _T_206 = _T_205 + _GEN_39; // @[GroupAllocator.scala 43:43:@13752.6]
  assign _T_207 = _T_205 + _GEN_39; // @[GroupAllocator.scala 43:43:@13753.6]
  assign _T_208 = io_storeHead - io_storeTail; // @[GroupAllocator.scala 45:22:@13757.6]
  assign _T_209 = $unsigned(_T_208); // @[GroupAllocator.scala 45:22:@13758.6]
  assign _T_210 = _T_209[2:0]; // @[GroupAllocator.scala 45:22:@13759.6]
  assign emptyStoreSlots = _T_201 ? _T_207 : {{1'd0}, _T_210}; // @[GroupAllocator.scala 42:34:@13748.4]
  assign _T_217 = 4'h1 <= emptyStoreSlots; // @[GroupAllocator.scala 54:19:@13765.4]
  assign _T_219 = 4'h2 <= emptyLoadSlots; // @[GroupAllocator.scala 54:50:@13766.4]
  assign possibleAllocations_0 = io_readyToPrevious_0 & io_bbStartSignals_0; // @[GroupAllocator.scala 56:106:@13773.4]
  assign possibleAllocations_1 = io_readyToPrevious_1 & io_bbStartSignals_1; // @[GroupAllocator.scala 56:106:@13774.4]
  assign allocatedBBIdx = possibleAllocations_0 ? 1'h0 : 1'h1; // @[Mux.scala 31:69:@13778.4]
  assign _T_244 = 1'h0 == allocatedBBIdx; // @[GroupAllocator.scala 69:43:@13782.4]
  assign _T_357 = allocatedBBIdx ? 2'h2 : 2'h0; // @[Mux.scala 46:16:@13872.6]
  assign _T_359 = _T_244 ? 2'h3 : _T_357; // @[Mux.scala 46:16:@13874.6]
  assign _T_368 = _T_244 ? 1'h0 : allocatedBBIdx; // @[Mux.scala 46:16:@13879.6]
  assign _T_438_0 = allocatedBBIdx ? 3'h3 : 3'h0; // @[Mux.scala 46:16:@13909.6]
  assign _T_438_1 = allocatedBBIdx ? 3'h4 : 3'h0; // @[Mux.scala 46:16:@13909.6]
  assign _T_459_0 = _T_244 ? 3'h0 : _T_438_0; // @[Mux.scala 46:16:@13911.6]
  assign _T_459_1 = _T_244 ? 3'h1 : _T_438_1; // @[Mux.scala 46:16:@13911.6]
  assign _T_459_2 = _T_244 ? 3'h2 : 3'h0; // @[Mux.scala 46:16:@13911.6]
  assign _T_614 = _GEN_38 + 4'h8; // @[GroupAllocator.scala 110:34:@13968.6]
  assign _T_615 = _GEN_38 + 4'h8; // @[GroupAllocator.scala 110:34:@13969.6]
  assign _T_617 = _T_615 - 4'h1; // @[GroupAllocator.scala 110:55:@13970.6]
  assign _T_618 = $unsigned(_T_617); // @[GroupAllocator.scala 110:55:@13971.6]
  assign _T_619 = _T_618[3:0]; // @[GroupAllocator.scala 110:55:@13972.6]
  assign _T_621 = {{1'd0}, _T_619}; // @[util.scala 10:8:@13973.6]
  assign _GEN_0 = _T_621 % 5'h8; // @[util.scala 10:14:@13974.6]
  assign _T_622 = _GEN_0[3:0]; // @[util.scala 10:14:@13974.6]
  assign _T_752 = _T_622[2:0]; // @[GroupAllocator.scala 110:90:@14056.6 GroupAllocator.scala 110:90:@14057.6]
  assign _T_866_0 = allocatedBBIdx ? _T_752 : 3'h0; // @[Mux.scala 46:16:@14131.6]
  assign _T_887_0 = _T_244 ? _T_752 : _T_866_0; // @[Mux.scala 46:16:@14133.6]
  assign _T_932 = _GEN_36 + 4'h8; // @[GroupAllocator.scala 115:33:@14151.6]
  assign _T_933 = _GEN_36 + 4'h8; // @[GroupAllocator.scala 115:33:@14152.6]
  assign _T_935 = _T_933 - 4'h1; // @[GroupAllocator.scala 115:54:@14153.6]
  assign _T_936 = $unsigned(_T_935); // @[GroupAllocator.scala 115:54:@14154.6]
  assign _T_937 = _T_936[3:0]; // @[GroupAllocator.scala 115:54:@14155.6]
  assign _T_939 = {{1'd0}, _T_937}; // @[util.scala 10:8:@14156.6]
  assign _GEN_1 = _T_939 % 5'h8; // @[util.scala 10:14:@14157.6]
  assign _T_940 = _GEN_1[3:0]; // @[util.scala 10:14:@14157.6]
  assign _T_1066 = 4'h2 + _T_937; // @[util.scala 10:8:@14237.6]
  assign _GEN_2 = _T_1066 % 5'h8; // @[util.scala 10:14:@14238.6]
  assign _T_1067 = _GEN_2[3:0]; // @[util.scala 10:14:@14238.6]
  assign _T_1070 = _T_1067[2:0]; // @[GroupAllocator.scala 115:89:@14239.6 GroupAllocator.scala 115:89:@14240.6]
  assign _T_1184_0 = allocatedBBIdx ? _T_1070 : 3'h0; // @[Mux.scala 46:16:@14314.6]
  assign _T_1084 = _T_940[2:0]; // @[GroupAllocator.scala 115:89:@14248.6 GroupAllocator.scala 115:89:@14249.6]
  assign _T_1184_1 = allocatedBBIdx ? _T_1084 : 3'h0; // @[Mux.scala 46:16:@14314.6]
  assign _T_1205_0 = _T_244 ? _T_1084 : _T_1184_0; // @[Mux.scala 46:16:@14316.6]
  assign _T_1205_1 = _T_244 ? _T_1084 : _T_1184_1; // @[Mux.scala 46:16:@14316.6]
  assign io_bbLoadOffsets_0 = io_bbStart ? _T_887_0 : 3'h0; // @[GroupAllocator.scala 89:20:@13845.4 GroupAllocator.scala 106:22:@14134.6]
  assign io_bbLoadOffsets_1 = io_bbStart ? _T_887_0 : 3'h0; // @[GroupAllocator.scala 89:20:@13846.4 GroupAllocator.scala 106:22:@14135.6]
  assign io_bbLoadOffsets_2 = io_bbStart ? _T_887_0 : 3'h0; // @[GroupAllocator.scala 89:20:@13847.4 GroupAllocator.scala 106:22:@14136.6]
  assign io_bbLoadOffsets_3 = io_bbStart ? _T_887_0 : 3'h0; // @[GroupAllocator.scala 89:20:@13848.4 GroupAllocator.scala 106:22:@14137.6]
  assign io_bbLoadOffsets_4 = io_bbStart ? _T_887_0 : 3'h0; // @[GroupAllocator.scala 89:20:@13849.4 GroupAllocator.scala 106:22:@14138.6]
  assign io_bbLoadOffsets_5 = io_bbStart ? _T_887_0 : 3'h0; // @[GroupAllocator.scala 89:20:@13850.4 GroupAllocator.scala 106:22:@14139.6]
  assign io_bbLoadOffsets_6 = io_bbStart ? _T_887_0 : 3'h0; // @[GroupAllocator.scala 89:20:@13851.4 GroupAllocator.scala 106:22:@14140.6]
  assign io_bbLoadOffsets_7 = io_bbStart ? _T_887_0 : 3'h0; // @[GroupAllocator.scala 89:20:@13852.4 GroupAllocator.scala 106:22:@14141.6]
  assign io_bbLoadPorts_0 = io_bbStart ? _T_459_0 : 3'h0; // @[GroupAllocator.scala 87:18:@13811.4 GroupAllocator.scala 95:20:@13912.6]
  assign io_bbLoadPorts_1 = io_bbStart ? _T_459_1 : 3'h0; // @[GroupAllocator.scala 87:18:@13812.4 GroupAllocator.scala 95:20:@13913.6]
  assign io_bbLoadPorts_2 = io_bbStart ? _T_459_2 : 3'h0; // @[GroupAllocator.scala 87:18:@13813.4 GroupAllocator.scala 95:20:@13914.6]
  assign io_bbNumLoads = io_bbStart ? {{1'd0}, _T_359} : 3'h0; // @[GroupAllocator.scala 85:17:@13800.4 GroupAllocator.scala 93:19:@13875.6]
  assign io_bbStoreOffsets_0 = io_bbStart ? _T_1205_0 : 3'h0; // @[GroupAllocator.scala 90:21:@13862.4 GroupAllocator.scala 111:23:@14317.6]
  assign io_bbStoreOffsets_1 = io_bbStart ? _T_1205_1 : 3'h0; // @[GroupAllocator.scala 90:21:@13863.4 GroupAllocator.scala 111:23:@14318.6]
  assign io_bbStoreOffsets_2 = io_bbStart ? _T_1205_1 : 3'h0; // @[GroupAllocator.scala 90:21:@13864.4 GroupAllocator.scala 111:23:@14319.6]
  assign io_bbStoreOffsets_3 = io_bbStart ? _T_1205_1 : 3'h0; // @[GroupAllocator.scala 90:21:@13865.4 GroupAllocator.scala 111:23:@14320.6]
  assign io_bbStoreOffsets_4 = io_bbStart ? _T_1205_1 : 3'h0; // @[GroupAllocator.scala 90:21:@13866.4 GroupAllocator.scala 111:23:@14321.6]
  assign io_bbStoreOffsets_5 = io_bbStart ? _T_1205_1 : 3'h0; // @[GroupAllocator.scala 90:21:@13867.4 GroupAllocator.scala 111:23:@14322.6]
  assign io_bbStoreOffsets_6 = io_bbStart ? _T_1205_1 : 3'h0; // @[GroupAllocator.scala 90:21:@13868.4 GroupAllocator.scala 111:23:@14323.6]
  assign io_bbStoreOffsets_7 = io_bbStart ? _T_1205_1 : 3'h0; // @[GroupAllocator.scala 90:21:@13869.4 GroupAllocator.scala 111:23:@14324.6]
  assign io_bbNumStores = io_bbStart ? _T_368 : 1'h0; // @[GroupAllocator.scala 86:18:@13801.4 GroupAllocator.scala 94:20:@13880.6]
  assign io_bbStart = possibleAllocations_0 | possibleAllocations_1; // @[GroupAllocator.scala 59:14:@13781.4]
  assign io_readyToPrevious_0 = 4'h3 <= emptyLoadSlots; // @[GroupAllocator.scala 53:22:@13771.4]
  assign io_readyToPrevious_1 = _T_217 & _T_219; // @[GroupAllocator.scala 53:22:@13772.4]
  assign io_loadPortsEnable_0 = _T_244 & io_bbStart; // @[GroupAllocator.scala 69:29:@13784.4]
  assign io_loadPortsEnable_1 = _T_244 & io_bbStart; // @[GroupAllocator.scala 69:29:@13787.4]
  assign io_loadPortsEnable_2 = _T_244 & io_bbStart; // @[GroupAllocator.scala 69:29:@13790.4]
  assign io_loadPortsEnable_3 = allocatedBBIdx & io_bbStart; // @[GroupAllocator.scala 69:29:@13793.4]
  assign io_loadPortsEnable_4 = allocatedBBIdx & io_bbStart; // @[GroupAllocator.scala 69:29:@13796.4]
  assign io_storePortsEnable_0 = allocatedBBIdx & io_bbStart; // @[GroupAllocator.scala 78:30:@13799.4]
endmodule
module LOAD_PORT_LSQ_dist( // @[:@14327.2]
  input         clock, // @[:@14328.4]
  input         reset, // @[:@14329.4]
  output        io_addrFromPrev_ready, // @[:@14330.4]
  input         io_addrFromPrev_valid, // @[:@14330.4]
  input  [31:0] io_addrFromPrev_bits, // @[:@14330.4]
  input         io_portEnable, // @[:@14330.4]
  input         io_dataToNext_ready, // @[:@14330.4]
  output        io_dataToNext_valid, // @[:@14330.4]
  output [31:0] io_dataToNext_bits, // @[:@14330.4]
  output        io_loadAddrEnable, // @[:@14330.4]
  output [31:0] io_addrToLoadQueue, // @[:@14330.4]
  output        io_dataFromLoadQueue_ready, // @[:@14330.4]
  input         io_dataFromLoadQueue_valid, // @[:@14330.4]
  input  [31:0] io_dataFromLoadQueue_bits // @[:@14330.4]
);
  reg [3:0] cnt; // @[LoadPort.scala 23:20:@14332.4]
  reg [31:0] _RAND_0;
  wire  _T_44; // @[LoadPort.scala 26:25:@14333.4]
  wire  _T_45; // @[LoadPort.scala 26:22:@14334.4]
  wire  _T_47; // @[LoadPort.scala 26:51:@14335.4]
  wire  _T_48; // @[LoadPort.scala 26:44:@14336.4]
  wire [4:0] _T_50; // @[LoadPort.scala 27:16:@14338.6]
  wire [3:0] _T_51; // @[LoadPort.scala 27:16:@14339.6]
  wire  _T_53; // @[LoadPort.scala 28:35:@14343.6]
  wire  _T_54; // @[LoadPort.scala 28:32:@14344.6]
  wire  _T_56; // @[LoadPort.scala 28:57:@14345.6]
  wire  _T_57; // @[LoadPort.scala 28:50:@14346.6]
  wire [4:0] _T_59; // @[LoadPort.scala 29:16:@14348.8]
  wire [4:0] _T_60; // @[LoadPort.scala 29:16:@14349.8]
  wire [3:0] _T_61; // @[LoadPort.scala 29:16:@14350.8]
  wire [3:0] _GEN_0; // @[LoadPort.scala 28:66:@14347.6]
  wire [3:0] _GEN_1; // @[LoadPort.scala 26:75:@14337.4]
  wire  _T_63; // @[LoadPort.scala 33:28:@14354.4]
  assign _T_44 = io_loadAddrEnable == 1'h0; // @[LoadPort.scala 26:25:@14333.4]
  assign _T_45 = io_portEnable & _T_44; // @[LoadPort.scala 26:22:@14334.4]
  assign _T_47 = cnt != 4'h8; // @[LoadPort.scala 26:51:@14335.4]
  assign _T_48 = _T_45 & _T_47; // @[LoadPort.scala 26:44:@14336.4]
  assign _T_50 = cnt + 4'h1; // @[LoadPort.scala 27:16:@14338.6]
  assign _T_51 = cnt + 4'h1; // @[LoadPort.scala 27:16:@14339.6]
  assign _T_53 = io_portEnable == 1'h0; // @[LoadPort.scala 28:35:@14343.6]
  assign _T_54 = io_loadAddrEnable & _T_53; // @[LoadPort.scala 28:32:@14344.6]
  assign _T_56 = cnt != 4'h0; // @[LoadPort.scala 28:57:@14345.6]
  assign _T_57 = _T_54 & _T_56; // @[LoadPort.scala 28:50:@14346.6]
  assign _T_59 = cnt - 4'h1; // @[LoadPort.scala 29:16:@14348.8]
  assign _T_60 = $unsigned(_T_59); // @[LoadPort.scala 29:16:@14349.8]
  assign _T_61 = _T_60[3:0]; // @[LoadPort.scala 29:16:@14350.8]
  assign _GEN_0 = _T_57 ? _T_61 : cnt; // @[LoadPort.scala 28:66:@14347.6]
  assign _GEN_1 = _T_48 ? _T_51 : _GEN_0; // @[LoadPort.scala 26:75:@14337.4]
  assign _T_63 = cnt > 4'h0; // @[LoadPort.scala 33:28:@14354.4]
  assign io_addrFromPrev_ready = cnt > 4'h0; // @[LoadPort.scala 34:25:@14358.4]
  assign io_dataToNext_valid = io_dataFromLoadQueue_valid; // @[LoadPort.scala 35:17:@14360.4]
  assign io_dataToNext_bits = io_dataFromLoadQueue_bits; // @[LoadPort.scala 35:17:@14359.4]
  assign io_loadAddrEnable = _T_63 & io_addrFromPrev_valid; // @[LoadPort.scala 33:21:@14356.4]
  assign io_addrToLoadQueue = io_addrFromPrev_bits; // @[LoadPort.scala 32:22:@14353.4]
  assign io_dataFromLoadQueue_ready = io_dataToNext_ready; // @[LoadPort.scala 35:17:@14361.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 4'h0;
    end else begin
      if (_T_48) begin
        cnt <= _T_51;
      end else begin
        if (_T_57) begin
          cnt <= _T_61;
        end
      end
    end
  end
endmodule
module STORE_DATA_PORT_LSQ_dist( // @[:@14507.2]
  input         clock, // @[:@14508.4]
  input         reset, // @[:@14509.4]
  output        io_dataFromPrev_ready, // @[:@14510.4]
  input         io_dataFromPrev_valid, // @[:@14510.4]
  input  [31:0] io_dataFromPrev_bits, // @[:@14510.4]
  input         io_portEnable, // @[:@14510.4]
  output        io_storeDataEnable, // @[:@14510.4]
  output [31:0] io_dataToStoreQueue // @[:@14510.4]
);
  reg [3:0] cnt; // @[StoreDataPort.scala 21:20:@14512.4]
  reg [31:0] _RAND_0;
  wire  _T_26; // @[StoreDataPort.scala 24:25:@14513.4]
  wire  _T_27; // @[StoreDataPort.scala 24:22:@14514.4]
  wire  _T_29; // @[StoreDataPort.scala 24:52:@14515.4]
  wire  _T_30; // @[StoreDataPort.scala 24:45:@14516.4]
  wire [4:0] _T_32; // @[StoreDataPort.scala 25:16:@14518.6]
  wire [3:0] _T_33; // @[StoreDataPort.scala 25:16:@14519.6]
  wire  _T_35; // @[StoreDataPort.scala 26:36:@14523.6]
  wire  _T_36; // @[StoreDataPort.scala 26:33:@14524.6]
  wire  _T_38; // @[StoreDataPort.scala 26:58:@14525.6]
  wire  _T_39; // @[StoreDataPort.scala 26:51:@14526.6]
  wire [4:0] _T_41; // @[StoreDataPort.scala 27:16:@14528.8]
  wire [4:0] _T_42; // @[StoreDataPort.scala 27:16:@14529.8]
  wire [3:0] _T_43; // @[StoreDataPort.scala 27:16:@14530.8]
  wire [3:0] _GEN_0; // @[StoreDataPort.scala 26:67:@14527.6]
  wire [3:0] _GEN_1; // @[StoreDataPort.scala 24:76:@14517.4]
  wire  _T_45; // @[StoreDataPort.scala 31:29:@14534.4]
  assign _T_26 = io_storeDataEnable == 1'h0; // @[StoreDataPort.scala 24:25:@14513.4]
  assign _T_27 = io_portEnable & _T_26; // @[StoreDataPort.scala 24:22:@14514.4]
  assign _T_29 = cnt != 4'h8; // @[StoreDataPort.scala 24:52:@14515.4]
  assign _T_30 = _T_27 & _T_29; // @[StoreDataPort.scala 24:45:@14516.4]
  assign _T_32 = cnt + 4'h1; // @[StoreDataPort.scala 25:16:@14518.6]
  assign _T_33 = cnt + 4'h1; // @[StoreDataPort.scala 25:16:@14519.6]
  assign _T_35 = io_portEnable == 1'h0; // @[StoreDataPort.scala 26:36:@14523.6]
  assign _T_36 = io_storeDataEnable & _T_35; // @[StoreDataPort.scala 26:33:@14524.6]
  assign _T_38 = cnt != 4'h0; // @[StoreDataPort.scala 26:58:@14525.6]
  assign _T_39 = _T_36 & _T_38; // @[StoreDataPort.scala 26:51:@14526.6]
  assign _T_41 = cnt - 4'h1; // @[StoreDataPort.scala 27:16:@14528.8]
  assign _T_42 = $unsigned(_T_41); // @[StoreDataPort.scala 27:16:@14529.8]
  assign _T_43 = _T_42[3:0]; // @[StoreDataPort.scala 27:16:@14530.8]
  assign _GEN_0 = _T_39 ? _T_43 : cnt; // @[StoreDataPort.scala 26:67:@14527.6]
  assign _GEN_1 = _T_30 ? _T_33 : _GEN_0; // @[StoreDataPort.scala 24:76:@14517.4]
  assign _T_45 = cnt > 4'h0; // @[StoreDataPort.scala 31:29:@14534.4]
  assign io_dataFromPrev_ready = cnt > 4'h0; // @[StoreDataPort.scala 32:25:@14538.4]
  assign io_storeDataEnable = _T_45 & io_dataFromPrev_valid; // @[StoreDataPort.scala 31:22:@14536.4]
  assign io_dataToStoreQueue = io_dataFromPrev_bits; // @[StoreDataPort.scala 30:23:@14533.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 4'h0;
    end else begin
      if (_T_30) begin
        cnt <= _T_33;
      end else begin
        if (_T_39) begin
          cnt <= _T_43;
        end
      end
    end
  end
endmodule
module LSQ_dist( // @[:@14573.2]
  input         clock, // @[:@14574.4]
  input         reset, // @[:@14575.4]
  output [31:0] io_storeDataOut, // @[:@14576.4]
  output [31:0] io_storeAddrOut, // @[:@14576.4]
  output        io_storeEnable, // @[:@14576.4]
  input         io_memIsReadyForStores, // @[:@14576.4]
  input  [31:0] io_loadDataIn, // @[:@14576.4]
  output [31:0] io_loadAddrOut, // @[:@14576.4]
  output        io_loadEnable, // @[:@14576.4]
  input         io_memIsReadyForLoads, // @[:@14576.4]
  input         io_bbpValids_0, // @[:@14576.4]
  input         io_bbpValids_1, // @[:@14576.4]
  output        io_bbReadyToPrevs_0, // @[:@14576.4]
  output        io_bbReadyToPrevs_1, // @[:@14576.4]
  output        io_rdPortsPrev_0_ready, // @[:@14576.4]
  input         io_rdPortsPrev_0_valid, // @[:@14576.4]
  input  [31:0] io_rdPortsPrev_0_bits, // @[:@14576.4]
  output        io_rdPortsPrev_1_ready, // @[:@14576.4]
  input         io_rdPortsPrev_1_valid, // @[:@14576.4]
  input  [31:0] io_rdPortsPrev_1_bits, // @[:@14576.4]
  output        io_rdPortsPrev_2_ready, // @[:@14576.4]
  input         io_rdPortsPrev_2_valid, // @[:@14576.4]
  input  [31:0] io_rdPortsPrev_2_bits, // @[:@14576.4]
  output        io_rdPortsPrev_3_ready, // @[:@14576.4]
  input         io_rdPortsPrev_3_valid, // @[:@14576.4]
  input  [31:0] io_rdPortsPrev_3_bits, // @[:@14576.4]
  output        io_rdPortsPrev_4_ready, // @[:@14576.4]
  input         io_rdPortsPrev_4_valid, // @[:@14576.4]
  input  [31:0] io_rdPortsPrev_4_bits, // @[:@14576.4]
  input         io_rdPortsNext_0_ready, // @[:@14576.4]
  output        io_rdPortsNext_0_valid, // @[:@14576.4]
  output [31:0] io_rdPortsNext_0_bits, // @[:@14576.4]
  input         io_rdPortsNext_1_ready, // @[:@14576.4]
  output        io_rdPortsNext_1_valid, // @[:@14576.4]
  output [31:0] io_rdPortsNext_1_bits, // @[:@14576.4]
  input         io_rdPortsNext_2_ready, // @[:@14576.4]
  output        io_rdPortsNext_2_valid, // @[:@14576.4]
  output [31:0] io_rdPortsNext_2_bits, // @[:@14576.4]
  input         io_rdPortsNext_3_ready, // @[:@14576.4]
  output        io_rdPortsNext_3_valid, // @[:@14576.4]
  output [31:0] io_rdPortsNext_3_bits, // @[:@14576.4]
  input         io_rdPortsNext_4_ready, // @[:@14576.4]
  output        io_rdPortsNext_4_valid, // @[:@14576.4]
  output [31:0] io_rdPortsNext_4_bits, // @[:@14576.4]
  output        io_wrAddrPorts_0_ready, // @[:@14576.4]
  input         io_wrAddrPorts_0_valid, // @[:@14576.4]
  input  [31:0] io_wrAddrPorts_0_bits, // @[:@14576.4]
  output        io_wrDataPorts_0_ready, // @[:@14576.4]
  input         io_wrDataPorts_0_valid, // @[:@14576.4]
  input  [31:0] io_wrDataPorts_0_bits, // @[:@14576.4]
  output        io_Empty_Valid // @[:@14576.4]
);
  wire  storeQ_clock; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_reset; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_bbStart; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_bbStoreOffsets_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_bbStoreOffsets_1; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_bbStoreOffsets_2; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_bbStoreOffsets_3; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_bbStoreOffsets_4; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_bbStoreOffsets_5; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_bbStoreOffsets_6; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_bbStoreOffsets_7; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_bbNumStores; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_storeTail; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_storeHead; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeEmpty; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_loadTail; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [2:0] storeQ_io_loadHead; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadEmpty; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadAddressDone_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadAddressDone_1; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadAddressDone_2; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadAddressDone_3; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadAddressDone_4; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadAddressDone_5; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadAddressDone_6; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadAddressDone_7; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadDataDone_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadDataDone_1; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadDataDone_2; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadDataDone_3; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadDataDone_4; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadDataDone_5; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadDataDone_6; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_loadDataDone_7; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_loadAddressQueue_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_loadAddressQueue_1; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_loadAddressQueue_2; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_loadAddressQueue_3; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_loadAddressQueue_4; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_loadAddressQueue_5; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_loadAddressQueue_6; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_loadAddressQueue_7; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeDataEnable_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_dataFromStorePorts_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeAddrEnable_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_addressFromStorePorts_0; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 72:22:@14607.4]
  wire [31:0] storeQ_io_storeDataToMem; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  storeQ_io_memIsReadyForStores; // @[LSQBRAM.scala 72:22:@14607.4]
  wire  loadQ_clock; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_reset; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_bbStart; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadOffsets_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadOffsets_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadOffsets_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadOffsets_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadOffsets_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadOffsets_5; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadOffsets_6; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadOffsets_7; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadPorts_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadPorts_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbLoadPorts_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_bbNumLoads; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_loadTail; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_loadHead; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadEmpty; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_storeTail; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] loadQ_io_storeHead; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeEmpty; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeAddrDone_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeAddrDone_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeAddrDone_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeAddrDone_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeAddrDone_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeAddrDone_5; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeAddrDone_6; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeAddrDone_7; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeDataDone_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeDataDone_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeDataDone_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeDataDone_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeDataDone_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeDataDone_5; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeDataDone_6; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_storeDataDone_7; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeDataQueue_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeDataQueue_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeDataQueue_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeDataQueue_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeDataQueue_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeDataQueue_5; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeDataQueue_6; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_storeDataQueue_7; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrEnable_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrEnable_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrEnable_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrEnable_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadAddrEnable_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_0; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_1; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_2; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_3; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_4; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_0_ready; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_1_ready; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_1_valid; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadPorts_1_bits; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_2_ready; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_2_valid; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadPorts_2_bits; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_3_ready; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_3_valid; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadPorts_3_bits; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_4_ready; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadPorts_4_valid; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadPorts_4_bits; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadDataFromMem; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [31:0] loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 73:21:@14610.4]
  wire  loadQ_io_memIsReadyForLoads; // @[LSQBRAM.scala 73:21:@14610.4]
  wire [2:0] GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadPorts_0; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadPorts_1; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbLoadPorts_2; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbNumLoads; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_loadTail; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_loadHead; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_loadEmpty; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_bbNumStores; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_storeTail; // @[LSQBRAM.scala 74:18:@14613.4]
  wire [2:0] GA_io_storeHead; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_storeEmpty; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_bbStart; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_bbStartSignals_0; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_bbStartSignals_1; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_readyToPrevious_0; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_readyToPrevious_1; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_loadPortsEnable_1; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_loadPortsEnable_2; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_loadPortsEnable_3; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_loadPortsEnable_4; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  GA_io_storePortsEnable_0; // @[LSQBRAM.scala 74:18:@14613.4]
  wire  LOAD_PORT_LSQ_dist_clock; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_reset; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@14616.4]
  wire [31:0] LOAD_PORT_LSQ_dist_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_io_portEnable; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@14616.4]
  wire [31:0] LOAD_PORT_LSQ_dist_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@14616.4]
  wire [31:0] LOAD_PORT_LSQ_dist_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@14616.4]
  wire [31:0] LOAD_PORT_LSQ_dist_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@14616.4]
  wire  LOAD_PORT_LSQ_dist_1_clock; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_1_reset; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_1_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_1_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@14619.4]
  wire [31:0] LOAD_PORT_LSQ_dist_1_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_1_io_portEnable; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_1_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_1_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@14619.4]
  wire [31:0] LOAD_PORT_LSQ_dist_1_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_1_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@14619.4]
  wire [31:0] LOAD_PORT_LSQ_dist_1_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_1_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_1_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@14619.4]
  wire [31:0] LOAD_PORT_LSQ_dist_1_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@14619.4]
  wire  LOAD_PORT_LSQ_dist_2_clock; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_2_reset; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_2_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_2_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@14622.4]
  wire [31:0] LOAD_PORT_LSQ_dist_2_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_2_io_portEnable; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_2_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_2_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@14622.4]
  wire [31:0] LOAD_PORT_LSQ_dist_2_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_2_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@14622.4]
  wire [31:0] LOAD_PORT_LSQ_dist_2_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_2_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_2_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@14622.4]
  wire [31:0] LOAD_PORT_LSQ_dist_2_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@14622.4]
  wire  LOAD_PORT_LSQ_dist_3_clock; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_3_reset; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_3_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_3_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@14625.4]
  wire [31:0] LOAD_PORT_LSQ_dist_3_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_3_io_portEnable; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_3_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_3_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@14625.4]
  wire [31:0] LOAD_PORT_LSQ_dist_3_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_3_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@14625.4]
  wire [31:0] LOAD_PORT_LSQ_dist_3_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_3_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_3_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@14625.4]
  wire [31:0] LOAD_PORT_LSQ_dist_3_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@14625.4]
  wire  LOAD_PORT_LSQ_dist_4_clock; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  LOAD_PORT_LSQ_dist_4_reset; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  LOAD_PORT_LSQ_dist_4_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  LOAD_PORT_LSQ_dist_4_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@14628.4]
  wire [31:0] LOAD_PORT_LSQ_dist_4_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  LOAD_PORT_LSQ_dist_4_io_portEnable; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  LOAD_PORT_LSQ_dist_4_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  LOAD_PORT_LSQ_dist_4_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@14628.4]
  wire [31:0] LOAD_PORT_LSQ_dist_4_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  LOAD_PORT_LSQ_dist_4_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@14628.4]
  wire [31:0] LOAD_PORT_LSQ_dist_4_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  LOAD_PORT_LSQ_dist_4_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  LOAD_PORT_LSQ_dist_4_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@14628.4]
  wire [31:0] LOAD_PORT_LSQ_dist_4_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@14628.4]
  wire  STORE_DATA_PORT_LSQ_dist_clock; // @[LSQBRAM.scala 80:11:@14692.4]
  wire  STORE_DATA_PORT_LSQ_dist_reset; // @[LSQBRAM.scala 80:11:@14692.4]
  wire  STORE_DATA_PORT_LSQ_dist_io_dataFromPrev_ready; // @[LSQBRAM.scala 80:11:@14692.4]
  wire  STORE_DATA_PORT_LSQ_dist_io_dataFromPrev_valid; // @[LSQBRAM.scala 80:11:@14692.4]
  wire [31:0] STORE_DATA_PORT_LSQ_dist_io_dataFromPrev_bits; // @[LSQBRAM.scala 80:11:@14692.4]
  wire  STORE_DATA_PORT_LSQ_dist_io_portEnable; // @[LSQBRAM.scala 80:11:@14692.4]
  wire  STORE_DATA_PORT_LSQ_dist_io_storeDataEnable; // @[LSQBRAM.scala 80:11:@14692.4]
  wire [31:0] STORE_DATA_PORT_LSQ_dist_io_dataToStoreQueue; // @[LSQBRAM.scala 80:11:@14692.4]
  wire  STORE_ADDR_PORT_LSQ_dist_clock; // @[LSQBRAM.scala 83:11:@14702.4]
  wire  STORE_ADDR_PORT_LSQ_dist_reset; // @[LSQBRAM.scala 83:11:@14702.4]
  wire  STORE_ADDR_PORT_LSQ_dist_io_dataFromPrev_ready; // @[LSQBRAM.scala 83:11:@14702.4]
  wire  STORE_ADDR_PORT_LSQ_dist_io_dataFromPrev_valid; // @[LSQBRAM.scala 83:11:@14702.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_dist_io_dataFromPrev_bits; // @[LSQBRAM.scala 83:11:@14702.4]
  wire  STORE_ADDR_PORT_LSQ_dist_io_portEnable; // @[LSQBRAM.scala 83:11:@14702.4]
  wire  STORE_ADDR_PORT_LSQ_dist_io_storeDataEnable; // @[LSQBRAM.scala 83:11:@14702.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_dist_io_dataToStoreQueue; // @[LSQBRAM.scala 83:11:@14702.4]
  wire  storeEmpty; // @[LSQBRAM.scala 46:24:@14583.4 LSQBRAM.scala 151:14:@14921.4]
  wire  loadEmpty; // @[LSQBRAM.scala 52:23:@14589.4 LSQBRAM.scala 119:13:@14820.4]
  wire [7:0] storeTail; // @[LSQBRAM.scala 44:23:@14581.4 LSQBRAM.scala 149:13:@14919.4]
  wire [7:0] storeHead; // @[LSQBRAM.scala 45:23:@14582.4 LSQBRAM.scala 150:13:@14920.4]
  wire [7:0] loadTail; // @[LSQBRAM.scala 50:22:@14587.4 LSQBRAM.scala 117:12:@14818.4]
  wire [7:0] loadHead; // @[LSQBRAM.scala 51:22:@14588.4 LSQBRAM.scala 118:12:@14819.4]
  STORE_QUEUE_LSQ_dist storeQ ( // @[LSQBRAM.scala 72:22:@14607.4]
    .clock(storeQ_clock),
    .reset(storeQ_reset),
    .io_bbStart(storeQ_io_bbStart),
    .io_bbStoreOffsets_0(storeQ_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(storeQ_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(storeQ_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(storeQ_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(storeQ_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(storeQ_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(storeQ_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(storeQ_io_bbStoreOffsets_7),
    .io_bbNumStores(storeQ_io_bbNumStores),
    .io_storeTail(storeQ_io_storeTail),
    .io_storeHead(storeQ_io_storeHead),
    .io_storeEmpty(storeQ_io_storeEmpty),
    .io_loadTail(storeQ_io_loadTail),
    .io_loadHead(storeQ_io_loadHead),
    .io_loadEmpty(storeQ_io_loadEmpty),
    .io_loadAddressDone_0(storeQ_io_loadAddressDone_0),
    .io_loadAddressDone_1(storeQ_io_loadAddressDone_1),
    .io_loadAddressDone_2(storeQ_io_loadAddressDone_2),
    .io_loadAddressDone_3(storeQ_io_loadAddressDone_3),
    .io_loadAddressDone_4(storeQ_io_loadAddressDone_4),
    .io_loadAddressDone_5(storeQ_io_loadAddressDone_5),
    .io_loadAddressDone_6(storeQ_io_loadAddressDone_6),
    .io_loadAddressDone_7(storeQ_io_loadAddressDone_7),
    .io_loadDataDone_0(storeQ_io_loadDataDone_0),
    .io_loadDataDone_1(storeQ_io_loadDataDone_1),
    .io_loadDataDone_2(storeQ_io_loadDataDone_2),
    .io_loadDataDone_3(storeQ_io_loadDataDone_3),
    .io_loadDataDone_4(storeQ_io_loadDataDone_4),
    .io_loadDataDone_5(storeQ_io_loadDataDone_5),
    .io_loadDataDone_6(storeQ_io_loadDataDone_6),
    .io_loadDataDone_7(storeQ_io_loadDataDone_7),
    .io_loadAddressQueue_0(storeQ_io_loadAddressQueue_0),
    .io_loadAddressQueue_1(storeQ_io_loadAddressQueue_1),
    .io_loadAddressQueue_2(storeQ_io_loadAddressQueue_2),
    .io_loadAddressQueue_3(storeQ_io_loadAddressQueue_3),
    .io_loadAddressQueue_4(storeQ_io_loadAddressQueue_4),
    .io_loadAddressQueue_5(storeQ_io_loadAddressQueue_5),
    .io_loadAddressQueue_6(storeQ_io_loadAddressQueue_6),
    .io_loadAddressQueue_7(storeQ_io_loadAddressQueue_7),
    .io_storeAddrDone_0(storeQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(storeQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(storeQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(storeQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(storeQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(storeQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(storeQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(storeQ_io_storeAddrDone_7),
    .io_storeDataDone_0(storeQ_io_storeDataDone_0),
    .io_storeDataDone_1(storeQ_io_storeDataDone_1),
    .io_storeDataDone_2(storeQ_io_storeDataDone_2),
    .io_storeDataDone_3(storeQ_io_storeDataDone_3),
    .io_storeDataDone_4(storeQ_io_storeDataDone_4),
    .io_storeDataDone_5(storeQ_io_storeDataDone_5),
    .io_storeDataDone_6(storeQ_io_storeDataDone_6),
    .io_storeDataDone_7(storeQ_io_storeDataDone_7),
    .io_storeAddrQueue_0(storeQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(storeQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(storeQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(storeQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(storeQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(storeQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(storeQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(storeQ_io_storeAddrQueue_7),
    .io_storeDataQueue_0(storeQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(storeQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(storeQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(storeQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(storeQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(storeQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(storeQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(storeQ_io_storeDataQueue_7),
    .io_storeDataEnable_0(storeQ_io_storeDataEnable_0),
    .io_dataFromStorePorts_0(storeQ_io_dataFromStorePorts_0),
    .io_storeAddrEnable_0(storeQ_io_storeAddrEnable_0),
    .io_addressFromStorePorts_0(storeQ_io_addressFromStorePorts_0),
    .io_storeAddrToMem(storeQ_io_storeAddrToMem),
    .io_storeDataToMem(storeQ_io_storeDataToMem),
    .io_storeEnableToMem(storeQ_io_storeEnableToMem),
    .io_memIsReadyForStores(storeQ_io_memIsReadyForStores)
  );
  LOAD_QUEUE_LSQ_dist loadQ ( // @[LSQBRAM.scala 73:21:@14610.4]
    .clock(loadQ_clock),
    .reset(loadQ_reset),
    .io_bbStart(loadQ_io_bbStart),
    .io_bbLoadOffsets_0(loadQ_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(loadQ_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(loadQ_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(loadQ_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(loadQ_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(loadQ_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(loadQ_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(loadQ_io_bbLoadOffsets_7),
    .io_bbLoadPorts_0(loadQ_io_bbLoadPorts_0),
    .io_bbLoadPorts_1(loadQ_io_bbLoadPorts_1),
    .io_bbLoadPorts_2(loadQ_io_bbLoadPorts_2),
    .io_bbNumLoads(loadQ_io_bbNumLoads),
    .io_loadTail(loadQ_io_loadTail),
    .io_loadHead(loadQ_io_loadHead),
    .io_loadEmpty(loadQ_io_loadEmpty),
    .io_storeTail(loadQ_io_storeTail),
    .io_storeHead(loadQ_io_storeHead),
    .io_storeEmpty(loadQ_io_storeEmpty),
    .io_storeAddrDone_0(loadQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(loadQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(loadQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(loadQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(loadQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(loadQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(loadQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(loadQ_io_storeAddrDone_7),
    .io_storeDataDone_0(loadQ_io_storeDataDone_0),
    .io_storeDataDone_1(loadQ_io_storeDataDone_1),
    .io_storeDataDone_2(loadQ_io_storeDataDone_2),
    .io_storeDataDone_3(loadQ_io_storeDataDone_3),
    .io_storeDataDone_4(loadQ_io_storeDataDone_4),
    .io_storeDataDone_5(loadQ_io_storeDataDone_5),
    .io_storeDataDone_6(loadQ_io_storeDataDone_6),
    .io_storeDataDone_7(loadQ_io_storeDataDone_7),
    .io_storeAddrQueue_0(loadQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(loadQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(loadQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(loadQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(loadQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(loadQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(loadQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(loadQ_io_storeAddrQueue_7),
    .io_storeDataQueue_0(loadQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(loadQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(loadQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(loadQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(loadQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(loadQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(loadQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(loadQ_io_storeDataQueue_7),
    .io_loadAddrDone_0(loadQ_io_loadAddrDone_0),
    .io_loadAddrDone_1(loadQ_io_loadAddrDone_1),
    .io_loadAddrDone_2(loadQ_io_loadAddrDone_2),
    .io_loadAddrDone_3(loadQ_io_loadAddrDone_3),
    .io_loadAddrDone_4(loadQ_io_loadAddrDone_4),
    .io_loadAddrDone_5(loadQ_io_loadAddrDone_5),
    .io_loadAddrDone_6(loadQ_io_loadAddrDone_6),
    .io_loadAddrDone_7(loadQ_io_loadAddrDone_7),
    .io_loadDataDone_0(loadQ_io_loadDataDone_0),
    .io_loadDataDone_1(loadQ_io_loadDataDone_1),
    .io_loadDataDone_2(loadQ_io_loadDataDone_2),
    .io_loadDataDone_3(loadQ_io_loadDataDone_3),
    .io_loadDataDone_4(loadQ_io_loadDataDone_4),
    .io_loadDataDone_5(loadQ_io_loadDataDone_5),
    .io_loadDataDone_6(loadQ_io_loadDataDone_6),
    .io_loadDataDone_7(loadQ_io_loadDataDone_7),
    .io_loadAddrQueue_0(loadQ_io_loadAddrQueue_0),
    .io_loadAddrQueue_1(loadQ_io_loadAddrQueue_1),
    .io_loadAddrQueue_2(loadQ_io_loadAddrQueue_2),
    .io_loadAddrQueue_3(loadQ_io_loadAddrQueue_3),
    .io_loadAddrQueue_4(loadQ_io_loadAddrQueue_4),
    .io_loadAddrQueue_5(loadQ_io_loadAddrQueue_5),
    .io_loadAddrQueue_6(loadQ_io_loadAddrQueue_6),
    .io_loadAddrQueue_7(loadQ_io_loadAddrQueue_7),
    .io_loadAddrEnable_0(loadQ_io_loadAddrEnable_0),
    .io_loadAddrEnable_1(loadQ_io_loadAddrEnable_1),
    .io_loadAddrEnable_2(loadQ_io_loadAddrEnable_2),
    .io_loadAddrEnable_3(loadQ_io_loadAddrEnable_3),
    .io_loadAddrEnable_4(loadQ_io_loadAddrEnable_4),
    .io_addrFromLoadPorts_0(loadQ_io_addrFromLoadPorts_0),
    .io_addrFromLoadPorts_1(loadQ_io_addrFromLoadPorts_1),
    .io_addrFromLoadPorts_2(loadQ_io_addrFromLoadPorts_2),
    .io_addrFromLoadPorts_3(loadQ_io_addrFromLoadPorts_3),
    .io_addrFromLoadPorts_4(loadQ_io_addrFromLoadPorts_4),
    .io_loadPorts_0_ready(loadQ_io_loadPorts_0_ready),
    .io_loadPorts_0_valid(loadQ_io_loadPorts_0_valid),
    .io_loadPorts_0_bits(loadQ_io_loadPorts_0_bits),
    .io_loadPorts_1_ready(loadQ_io_loadPorts_1_ready),
    .io_loadPorts_1_valid(loadQ_io_loadPorts_1_valid),
    .io_loadPorts_1_bits(loadQ_io_loadPorts_1_bits),
    .io_loadPorts_2_ready(loadQ_io_loadPorts_2_ready),
    .io_loadPorts_2_valid(loadQ_io_loadPorts_2_valid),
    .io_loadPorts_2_bits(loadQ_io_loadPorts_2_bits),
    .io_loadPorts_3_ready(loadQ_io_loadPorts_3_ready),
    .io_loadPorts_3_valid(loadQ_io_loadPorts_3_valid),
    .io_loadPorts_3_bits(loadQ_io_loadPorts_3_bits),
    .io_loadPorts_4_ready(loadQ_io_loadPorts_4_ready),
    .io_loadPorts_4_valid(loadQ_io_loadPorts_4_valid),
    .io_loadPorts_4_bits(loadQ_io_loadPorts_4_bits),
    .io_loadDataFromMem(loadQ_io_loadDataFromMem),
    .io_loadAddrToMem(loadQ_io_loadAddrToMem),
    .io_loadEnableToMem(loadQ_io_loadEnableToMem),
    .io_memIsReadyForLoads(loadQ_io_memIsReadyForLoads)
  );
  GROUP_ALLOCATOR_LSQ_dist GA ( // @[LSQBRAM.scala 74:18:@14613.4]
    .io_bbLoadOffsets_0(GA_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(GA_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(GA_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(GA_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(GA_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(GA_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(GA_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(GA_io_bbLoadOffsets_7),
    .io_bbLoadPorts_0(GA_io_bbLoadPorts_0),
    .io_bbLoadPorts_1(GA_io_bbLoadPorts_1),
    .io_bbLoadPorts_2(GA_io_bbLoadPorts_2),
    .io_bbNumLoads(GA_io_bbNumLoads),
    .io_loadTail(GA_io_loadTail),
    .io_loadHead(GA_io_loadHead),
    .io_loadEmpty(GA_io_loadEmpty),
    .io_bbStoreOffsets_0(GA_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(GA_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(GA_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(GA_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(GA_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(GA_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(GA_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(GA_io_bbStoreOffsets_7),
    .io_bbNumStores(GA_io_bbNumStores),
    .io_storeTail(GA_io_storeTail),
    .io_storeHead(GA_io_storeHead),
    .io_storeEmpty(GA_io_storeEmpty),
    .io_bbStart(GA_io_bbStart),
    .io_bbStartSignals_0(GA_io_bbStartSignals_0),
    .io_bbStartSignals_1(GA_io_bbStartSignals_1),
    .io_readyToPrevious_0(GA_io_readyToPrevious_0),
    .io_readyToPrevious_1(GA_io_readyToPrevious_1),
    .io_loadPortsEnable_0(GA_io_loadPortsEnable_0),
    .io_loadPortsEnable_1(GA_io_loadPortsEnable_1),
    .io_loadPortsEnable_2(GA_io_loadPortsEnable_2),
    .io_loadPortsEnable_3(GA_io_loadPortsEnable_3),
    .io_loadPortsEnable_4(GA_io_loadPortsEnable_4),
    .io_storePortsEnable_0(GA_io_storePortsEnable_0)
  );
  LOAD_PORT_LSQ_dist LOAD_PORT_LSQ_dist ( // @[LSQBRAM.scala 77:11:@14616.4]
    .clock(LOAD_PORT_LSQ_dist_clock),
    .reset(LOAD_PORT_LSQ_dist_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_dist_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_dist_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_dist_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_dist_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_dist_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_dist_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_dist_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_dist_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_dist_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_dist_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_dist_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_dist_io_dataFromLoadQueue_bits)
  );
  LOAD_PORT_LSQ_dist LOAD_PORT_LSQ_dist_1 ( // @[LSQBRAM.scala 77:11:@14619.4]
    .clock(LOAD_PORT_LSQ_dist_1_clock),
    .reset(LOAD_PORT_LSQ_dist_1_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_dist_1_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_dist_1_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_dist_1_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_dist_1_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_dist_1_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_dist_1_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_dist_1_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_dist_1_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_dist_1_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_dist_1_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_dist_1_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_dist_1_io_dataFromLoadQueue_bits)
  );
  LOAD_PORT_LSQ_dist LOAD_PORT_LSQ_dist_2 ( // @[LSQBRAM.scala 77:11:@14622.4]
    .clock(LOAD_PORT_LSQ_dist_2_clock),
    .reset(LOAD_PORT_LSQ_dist_2_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_dist_2_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_dist_2_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_dist_2_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_dist_2_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_dist_2_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_dist_2_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_dist_2_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_dist_2_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_dist_2_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_dist_2_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_dist_2_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_dist_2_io_dataFromLoadQueue_bits)
  );
  LOAD_PORT_LSQ_dist LOAD_PORT_LSQ_dist_3 ( // @[LSQBRAM.scala 77:11:@14625.4]
    .clock(LOAD_PORT_LSQ_dist_3_clock),
    .reset(LOAD_PORT_LSQ_dist_3_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_dist_3_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_dist_3_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_dist_3_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_dist_3_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_dist_3_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_dist_3_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_dist_3_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_dist_3_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_dist_3_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_dist_3_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_dist_3_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_dist_3_io_dataFromLoadQueue_bits)
  );
  LOAD_PORT_LSQ_dist LOAD_PORT_LSQ_dist_4 ( // @[LSQBRAM.scala 77:11:@14628.4]
    .clock(LOAD_PORT_LSQ_dist_4_clock),
    .reset(LOAD_PORT_LSQ_dist_4_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_dist_4_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_dist_4_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_dist_4_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_dist_4_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_dist_4_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_dist_4_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_dist_4_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_dist_4_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_dist_4_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_dist_4_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_dist_4_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_dist_4_io_dataFromLoadQueue_bits)
  );
  STORE_DATA_PORT_LSQ_dist STORE_DATA_PORT_LSQ_dist ( // @[LSQBRAM.scala 80:11:@14692.4]
    .clock(STORE_DATA_PORT_LSQ_dist_clock),
    .reset(STORE_DATA_PORT_LSQ_dist_reset),
    .io_dataFromPrev_ready(STORE_DATA_PORT_LSQ_dist_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_DATA_PORT_LSQ_dist_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_DATA_PORT_LSQ_dist_io_dataFromPrev_bits),
    .io_portEnable(STORE_DATA_PORT_LSQ_dist_io_portEnable),
    .io_storeDataEnable(STORE_DATA_PORT_LSQ_dist_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_DATA_PORT_LSQ_dist_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_dist STORE_ADDR_PORT_LSQ_dist ( // @[LSQBRAM.scala 83:11:@14702.4]
    .clock(STORE_ADDR_PORT_LSQ_dist_clock),
    .reset(STORE_ADDR_PORT_LSQ_dist_reset),
    .io_dataFromPrev_ready(STORE_ADDR_PORT_LSQ_dist_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_ADDR_PORT_LSQ_dist_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_ADDR_PORT_LSQ_dist_io_dataFromPrev_bits),
    .io_portEnable(STORE_ADDR_PORT_LSQ_dist_io_portEnable),
    .io_storeDataEnable(STORE_ADDR_PORT_LSQ_dist_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_ADDR_PORT_LSQ_dist_io_dataToStoreQueue)
  );
  assign storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 46:24:@14583.4 LSQBRAM.scala 151:14:@14921.4]
  assign loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 52:23:@14589.4 LSQBRAM.scala 119:13:@14820.4]
  assign storeTail = {{5'd0}, storeQ_io_storeTail}; // @[LSQBRAM.scala 44:23:@14581.4 LSQBRAM.scala 149:13:@14919.4]
  assign storeHead = {{5'd0}, storeQ_io_storeHead}; // @[LSQBRAM.scala 45:23:@14582.4 LSQBRAM.scala 150:13:@14920.4]
  assign loadTail = {{5'd0}, loadQ_io_loadTail}; // @[LSQBRAM.scala 50:22:@14587.4 LSQBRAM.scala 117:12:@14818.4]
  assign loadHead = {{5'd0}, loadQ_io_loadHead}; // @[LSQBRAM.scala 51:22:@14588.4 LSQBRAM.scala 118:12:@14819.4]
  assign io_storeDataOut = storeQ_io_storeDataToMem; // @[LSQBRAM.scala 161:19:@14959.4]
  assign io_storeAddrOut = storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 160:19:@14958.4]
  assign io_storeEnable = storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 162:18:@14960.4]
  assign io_loadAddrOut = loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 135:18:@14872.4]
  assign io_loadEnable = loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 136:17:@14873.4]
  assign io_bbReadyToPrevs_0 = GA_io_readyToPrevious_0; // @[LSQBRAM.scala 102:21:@14757.4]
  assign io_bbReadyToPrevs_1 = GA_io_readyToPrevious_1; // @[LSQBRAM.scala 102:21:@14758.4]
  assign io_rdPortsPrev_0_ready = LOAD_PORT_LSQ_dist_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@14964.4]
  assign io_rdPortsPrev_1_ready = LOAD_PORT_LSQ_dist_1_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@14976.4]
  assign io_rdPortsPrev_2_ready = LOAD_PORT_LSQ_dist_2_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@14988.4]
  assign io_rdPortsPrev_3_ready = LOAD_PORT_LSQ_dist_3_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@15000.4]
  assign io_rdPortsPrev_4_ready = LOAD_PORT_LSQ_dist_4_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@15012.4]
  assign io_rdPortsNext_0_valid = LOAD_PORT_LSQ_dist_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@14967.4]
  assign io_rdPortsNext_0_bits = LOAD_PORT_LSQ_dist_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@14966.4]
  assign io_rdPortsNext_1_valid = LOAD_PORT_LSQ_dist_1_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@14979.4]
  assign io_rdPortsNext_1_bits = LOAD_PORT_LSQ_dist_1_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@14978.4]
  assign io_rdPortsNext_2_valid = LOAD_PORT_LSQ_dist_2_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@14991.4]
  assign io_rdPortsNext_2_bits = LOAD_PORT_LSQ_dist_2_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@14990.4]
  assign io_rdPortsNext_3_valid = LOAD_PORT_LSQ_dist_3_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@15003.4]
  assign io_rdPortsNext_3_bits = LOAD_PORT_LSQ_dist_3_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@15002.4]
  assign io_rdPortsNext_4_valid = LOAD_PORT_LSQ_dist_4_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@15015.4]
  assign io_rdPortsNext_4_bits = LOAD_PORT_LSQ_dist_4_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@15014.4]
  assign io_wrAddrPorts_0_ready = STORE_ADDR_PORT_LSQ_dist_io_dataFromPrev_ready; // @[LSQBRAM.scala 182:39:@15030.4]
  assign io_wrDataPorts_0_ready = STORE_DATA_PORT_LSQ_dist_io_dataFromPrev_ready; // @[LSQBRAM.scala 177:36:@15024.4]
  assign io_Empty_Valid = storeEmpty & loadEmpty; // @[LSQBRAM.scala 86:18:@14713.4]
  assign storeQ_clock = clock; // @[:@14608.4]
  assign storeQ_reset = reset; // @[:@14609.4]
  assign storeQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 145:21:@14901.4]
  assign storeQ_io_bbStoreOffsets_0 = GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 146:28:@14902.4]
  assign storeQ_io_bbStoreOffsets_1 = GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 146:28:@14903.4]
  assign storeQ_io_bbStoreOffsets_2 = GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 146:28:@14904.4]
  assign storeQ_io_bbStoreOffsets_3 = GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 146:28:@14905.4]
  assign storeQ_io_bbStoreOffsets_4 = GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 146:28:@14906.4]
  assign storeQ_io_bbStoreOffsets_5 = GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 146:28:@14907.4]
  assign storeQ_io_bbStoreOffsets_6 = GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 146:28:@14908.4]
  assign storeQ_io_bbStoreOffsets_7 = GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 146:28:@14909.4]
  assign storeQ_io_bbNumStores = {{2'd0}, GA_io_bbNumStores}; // @[LSQBRAM.scala 148:25:@14918.4]
  assign storeQ_io_loadTail = loadTail[2:0]; // @[LSQBRAM.scala 139:22:@14874.4]
  assign storeQ_io_loadHead = loadHead[2:0]; // @[LSQBRAM.scala 140:22:@14875.4]
  assign storeQ_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 141:23:@14876.4]
  assign storeQ_io_loadAddressDone_0 = loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 142:29:@14877.4]
  assign storeQ_io_loadAddressDone_1 = loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 142:29:@14878.4]
  assign storeQ_io_loadAddressDone_2 = loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 142:29:@14879.4]
  assign storeQ_io_loadAddressDone_3 = loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 142:29:@14880.4]
  assign storeQ_io_loadAddressDone_4 = loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 142:29:@14881.4]
  assign storeQ_io_loadAddressDone_5 = loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 142:29:@14882.4]
  assign storeQ_io_loadAddressDone_6 = loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 142:29:@14883.4]
  assign storeQ_io_loadAddressDone_7 = loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 142:29:@14884.4]
  assign storeQ_io_loadDataDone_0 = loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 143:26:@14885.4]
  assign storeQ_io_loadDataDone_1 = loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 143:26:@14886.4]
  assign storeQ_io_loadDataDone_2 = loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 143:26:@14887.4]
  assign storeQ_io_loadDataDone_3 = loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 143:26:@14888.4]
  assign storeQ_io_loadDataDone_4 = loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 143:26:@14889.4]
  assign storeQ_io_loadDataDone_5 = loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 143:26:@14890.4]
  assign storeQ_io_loadDataDone_6 = loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 143:26:@14891.4]
  assign storeQ_io_loadDataDone_7 = loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 143:26:@14892.4]
  assign storeQ_io_loadAddressQueue_0 = loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 144:30:@14893.4]
  assign storeQ_io_loadAddressQueue_1 = loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 144:30:@14894.4]
  assign storeQ_io_loadAddressQueue_2 = loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 144:30:@14895.4]
  assign storeQ_io_loadAddressQueue_3 = loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 144:30:@14896.4]
  assign storeQ_io_loadAddressQueue_4 = loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 144:30:@14897.4]
  assign storeQ_io_loadAddressQueue_5 = loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 144:30:@14898.4]
  assign storeQ_io_loadAddressQueue_6 = loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 144:30:@14899.4]
  assign storeQ_io_loadAddressQueue_7 = loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 144:30:@14900.4]
  assign storeQ_io_storeDataEnable_0 = STORE_DATA_PORT_LSQ_dist_io_storeDataEnable; // @[LSQBRAM.scala 156:29:@14954.4]
  assign storeQ_io_dataFromStorePorts_0 = STORE_DATA_PORT_LSQ_dist_io_dataToStoreQueue; // @[LSQBRAM.scala 157:32:@14955.4]
  assign storeQ_io_storeAddrEnable_0 = STORE_ADDR_PORT_LSQ_dist_io_storeDataEnable; // @[LSQBRAM.scala 158:29:@14956.4]
  assign storeQ_io_addressFromStorePorts_0 = STORE_ADDR_PORT_LSQ_dist_io_dataToStoreQueue; // @[LSQBRAM.scala 159:35:@14957.4]
  assign storeQ_io_memIsReadyForStores = io_memIsReadyForStores; // @[LSQBRAM.scala 163:33:@14961.4]
  assign loadQ_clock = clock; // @[:@14611.4]
  assign loadQ_reset = reset; // @[:@14612.4]
  assign loadQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 113:20:@14800.4]
  assign loadQ_io_bbLoadOffsets_0 = GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 114:26:@14801.4]
  assign loadQ_io_bbLoadOffsets_1 = GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 114:26:@14802.4]
  assign loadQ_io_bbLoadOffsets_2 = GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 114:26:@14803.4]
  assign loadQ_io_bbLoadOffsets_3 = GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 114:26:@14804.4]
  assign loadQ_io_bbLoadOffsets_4 = GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 114:26:@14805.4]
  assign loadQ_io_bbLoadOffsets_5 = GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 114:26:@14806.4]
  assign loadQ_io_bbLoadOffsets_6 = GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 114:26:@14807.4]
  assign loadQ_io_bbLoadOffsets_7 = GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 114:26:@14808.4]
  assign loadQ_io_bbLoadPorts_0 = GA_io_bbLoadPorts_0; // @[LSQBRAM.scala 115:24:@14809.4]
  assign loadQ_io_bbLoadPorts_1 = GA_io_bbLoadPorts_1; // @[LSQBRAM.scala 115:24:@14810.4]
  assign loadQ_io_bbLoadPorts_2 = GA_io_bbLoadPorts_2; // @[LSQBRAM.scala 115:24:@14811.4]
  assign loadQ_io_bbNumLoads = GA_io_bbNumLoads; // @[LSQBRAM.scala 116:23:@14817.4]
  assign loadQ_io_storeTail = storeTail[2:0]; // @[LSQBRAM.scala 106:22:@14765.4]
  assign loadQ_io_storeHead = storeHead[2:0]; // @[LSQBRAM.scala 107:22:@14766.4]
  assign loadQ_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 108:23:@14767.4]
  assign loadQ_io_storeAddrDone_0 = storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 109:26:@14768.4]
  assign loadQ_io_storeAddrDone_1 = storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 109:26:@14769.4]
  assign loadQ_io_storeAddrDone_2 = storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 109:26:@14770.4]
  assign loadQ_io_storeAddrDone_3 = storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 109:26:@14771.4]
  assign loadQ_io_storeAddrDone_4 = storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 109:26:@14772.4]
  assign loadQ_io_storeAddrDone_5 = storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 109:26:@14773.4]
  assign loadQ_io_storeAddrDone_6 = storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 109:26:@14774.4]
  assign loadQ_io_storeAddrDone_7 = storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 109:26:@14775.4]
  assign loadQ_io_storeDataDone_0 = storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 110:26:@14776.4]
  assign loadQ_io_storeDataDone_1 = storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 110:26:@14777.4]
  assign loadQ_io_storeDataDone_2 = storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 110:26:@14778.4]
  assign loadQ_io_storeDataDone_3 = storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 110:26:@14779.4]
  assign loadQ_io_storeDataDone_4 = storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 110:26:@14780.4]
  assign loadQ_io_storeDataDone_5 = storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 110:26:@14781.4]
  assign loadQ_io_storeDataDone_6 = storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 110:26:@14782.4]
  assign loadQ_io_storeDataDone_7 = storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 110:26:@14783.4]
  assign loadQ_io_storeAddrQueue_0 = storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 111:27:@14784.4]
  assign loadQ_io_storeAddrQueue_1 = storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 111:27:@14785.4]
  assign loadQ_io_storeAddrQueue_2 = storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 111:27:@14786.4]
  assign loadQ_io_storeAddrQueue_3 = storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 111:27:@14787.4]
  assign loadQ_io_storeAddrQueue_4 = storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 111:27:@14788.4]
  assign loadQ_io_storeAddrQueue_5 = storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 111:27:@14789.4]
  assign loadQ_io_storeAddrQueue_6 = storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 111:27:@14790.4]
  assign loadQ_io_storeAddrQueue_7 = storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 111:27:@14791.4]
  assign loadQ_io_storeDataQueue_0 = storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 112:27:@14792.4]
  assign loadQ_io_storeDataQueue_1 = storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 112:27:@14793.4]
  assign loadQ_io_storeDataQueue_2 = storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 112:27:@14794.4]
  assign loadQ_io_storeDataQueue_3 = storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 112:27:@14795.4]
  assign loadQ_io_storeDataQueue_4 = storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 112:27:@14796.4]
  assign loadQ_io_storeDataQueue_5 = storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 112:27:@14797.4]
  assign loadQ_io_storeDataQueue_6 = storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 112:27:@14798.4]
  assign loadQ_io_storeDataQueue_7 = storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 112:27:@14799.4]
  assign loadQ_io_loadAddrEnable_0 = LOAD_PORT_LSQ_dist_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@14849.4]
  assign loadQ_io_loadAddrEnable_1 = LOAD_PORT_LSQ_dist_1_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@14854.4]
  assign loadQ_io_loadAddrEnable_2 = LOAD_PORT_LSQ_dist_2_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@14859.4]
  assign loadQ_io_loadAddrEnable_3 = LOAD_PORT_LSQ_dist_3_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@14864.4]
  assign loadQ_io_loadAddrEnable_4 = LOAD_PORT_LSQ_dist_4_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@14869.4]
  assign loadQ_io_addrFromLoadPorts_0 = LOAD_PORT_LSQ_dist_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@14848.4]
  assign loadQ_io_addrFromLoadPorts_1 = LOAD_PORT_LSQ_dist_1_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@14853.4]
  assign loadQ_io_addrFromLoadPorts_2 = LOAD_PORT_LSQ_dist_2_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@14858.4]
  assign loadQ_io_addrFromLoadPorts_3 = LOAD_PORT_LSQ_dist_3_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@14863.4]
  assign loadQ_io_addrFromLoadPorts_4 = LOAD_PORT_LSQ_dist_4_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@14868.4]
  assign loadQ_io_loadPorts_0_ready = LOAD_PORT_LSQ_dist_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@14847.4]
  assign loadQ_io_loadPorts_1_ready = LOAD_PORT_LSQ_dist_1_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@14852.4]
  assign loadQ_io_loadPorts_2_ready = LOAD_PORT_LSQ_dist_2_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@14857.4]
  assign loadQ_io_loadPorts_3_ready = LOAD_PORT_LSQ_dist_3_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@14862.4]
  assign loadQ_io_loadPorts_4_ready = LOAD_PORT_LSQ_dist_4_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@14867.4]
  assign loadQ_io_loadDataFromMem = io_loadDataIn; // @[LSQBRAM.scala 133:28:@14870.4]
  assign loadQ_io_memIsReadyForLoads = io_memIsReadyForLoads; // @[LSQBRAM.scala 134:31:@14871.4]
  assign GA_io_loadTail = loadTail[2:0]; // @[LSQBRAM.scala 91:18:@14731.4]
  assign GA_io_loadHead = loadHead[2:0]; // @[LSQBRAM.scala 92:18:@14732.4]
  assign GA_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 93:19:@14733.4]
  assign GA_io_storeTail = storeTail[2:0]; // @[LSQBRAM.scala 97:19:@14751.4]
  assign GA_io_storeHead = storeHead[2:0]; // @[LSQBRAM.scala 98:19:@14752.4]
  assign GA_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 99:20:@14753.4]
  assign GA_io_bbStartSignals_0 = io_bbpValids_0; // @[LSQBRAM.scala 101:24:@14755.4]
  assign GA_io_bbStartSignals_1 = io_bbpValids_1; // @[LSQBRAM.scala 101:24:@14756.4]
  assign LOAD_PORT_LSQ_dist_clock = clock; // @[:@14617.4]
  assign LOAD_PORT_LSQ_dist_reset = reset; // @[:@14618.4]
  assign LOAD_PORT_LSQ_dist_io_addrFromPrev_valid = io_rdPortsPrev_0_valid; // @[LSQBRAM.scala 76:26:@14642.4]
  assign LOAD_PORT_LSQ_dist_io_addrFromPrev_bits = io_rdPortsPrev_0_bits; // @[LSQBRAM.scala 76:26:@14641.4]
  assign LOAD_PORT_LSQ_dist_io_portEnable = GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 76:26:@14640.4]
  assign LOAD_PORT_LSQ_dist_io_dataToNext_ready = io_rdPortsNext_0_ready; // @[LSQBRAM.scala 76:26:@14639.4]
  assign LOAD_PORT_LSQ_dist_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 76:26:@14633.4]
  assign LOAD_PORT_LSQ_dist_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 76:26:@14632.4]
  assign LOAD_PORT_LSQ_dist_1_clock = clock; // @[:@14620.4]
  assign LOAD_PORT_LSQ_dist_1_reset = reset; // @[:@14621.4]
  assign LOAD_PORT_LSQ_dist_1_io_addrFromPrev_valid = io_rdPortsPrev_1_valid; // @[LSQBRAM.scala 76:26:@14654.4]
  assign LOAD_PORT_LSQ_dist_1_io_addrFromPrev_bits = io_rdPortsPrev_1_bits; // @[LSQBRAM.scala 76:26:@14653.4]
  assign LOAD_PORT_LSQ_dist_1_io_portEnable = GA_io_loadPortsEnable_1; // @[LSQBRAM.scala 76:26:@14652.4]
  assign LOAD_PORT_LSQ_dist_1_io_dataToNext_ready = io_rdPortsNext_1_ready; // @[LSQBRAM.scala 76:26:@14651.4]
  assign LOAD_PORT_LSQ_dist_1_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_1_valid; // @[LSQBRAM.scala 76:26:@14645.4]
  assign LOAD_PORT_LSQ_dist_1_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_1_bits; // @[LSQBRAM.scala 76:26:@14644.4]
  assign LOAD_PORT_LSQ_dist_2_clock = clock; // @[:@14623.4]
  assign LOAD_PORT_LSQ_dist_2_reset = reset; // @[:@14624.4]
  assign LOAD_PORT_LSQ_dist_2_io_addrFromPrev_valid = io_rdPortsPrev_2_valid; // @[LSQBRAM.scala 76:26:@14666.4]
  assign LOAD_PORT_LSQ_dist_2_io_addrFromPrev_bits = io_rdPortsPrev_2_bits; // @[LSQBRAM.scala 76:26:@14665.4]
  assign LOAD_PORT_LSQ_dist_2_io_portEnable = GA_io_loadPortsEnable_2; // @[LSQBRAM.scala 76:26:@14664.4]
  assign LOAD_PORT_LSQ_dist_2_io_dataToNext_ready = io_rdPortsNext_2_ready; // @[LSQBRAM.scala 76:26:@14663.4]
  assign LOAD_PORT_LSQ_dist_2_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_2_valid; // @[LSQBRAM.scala 76:26:@14657.4]
  assign LOAD_PORT_LSQ_dist_2_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_2_bits; // @[LSQBRAM.scala 76:26:@14656.4]
  assign LOAD_PORT_LSQ_dist_3_clock = clock; // @[:@14626.4]
  assign LOAD_PORT_LSQ_dist_3_reset = reset; // @[:@14627.4]
  assign LOAD_PORT_LSQ_dist_3_io_addrFromPrev_valid = io_rdPortsPrev_3_valid; // @[LSQBRAM.scala 76:26:@14678.4]
  assign LOAD_PORT_LSQ_dist_3_io_addrFromPrev_bits = io_rdPortsPrev_3_bits; // @[LSQBRAM.scala 76:26:@14677.4]
  assign LOAD_PORT_LSQ_dist_3_io_portEnable = GA_io_loadPortsEnable_3; // @[LSQBRAM.scala 76:26:@14676.4]
  assign LOAD_PORT_LSQ_dist_3_io_dataToNext_ready = io_rdPortsNext_3_ready; // @[LSQBRAM.scala 76:26:@14675.4]
  assign LOAD_PORT_LSQ_dist_3_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_3_valid; // @[LSQBRAM.scala 76:26:@14669.4]
  assign LOAD_PORT_LSQ_dist_3_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_3_bits; // @[LSQBRAM.scala 76:26:@14668.4]
  assign LOAD_PORT_LSQ_dist_4_clock = clock; // @[:@14629.4]
  assign LOAD_PORT_LSQ_dist_4_reset = reset; // @[:@14630.4]
  assign LOAD_PORT_LSQ_dist_4_io_addrFromPrev_valid = io_rdPortsPrev_4_valid; // @[LSQBRAM.scala 76:26:@14690.4]
  assign LOAD_PORT_LSQ_dist_4_io_addrFromPrev_bits = io_rdPortsPrev_4_bits; // @[LSQBRAM.scala 76:26:@14689.4]
  assign LOAD_PORT_LSQ_dist_4_io_portEnable = GA_io_loadPortsEnable_4; // @[LSQBRAM.scala 76:26:@14688.4]
  assign LOAD_PORT_LSQ_dist_4_io_dataToNext_ready = io_rdPortsNext_4_ready; // @[LSQBRAM.scala 76:26:@14687.4]
  assign LOAD_PORT_LSQ_dist_4_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_4_valid; // @[LSQBRAM.scala 76:26:@14681.4]
  assign LOAD_PORT_LSQ_dist_4_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_4_bits; // @[LSQBRAM.scala 76:26:@14680.4]
  assign STORE_DATA_PORT_LSQ_dist_clock = clock; // @[:@14693.4]
  assign STORE_DATA_PORT_LSQ_dist_reset = reset; // @[:@14694.4]
  assign STORE_DATA_PORT_LSQ_dist_io_dataFromPrev_valid = io_wrDataPorts_0_valid; // @[LSQBRAM.scala 79:31:@14700.4]
  assign STORE_DATA_PORT_LSQ_dist_io_dataFromPrev_bits = io_wrDataPorts_0_bits; // @[LSQBRAM.scala 79:31:@14699.4]
  assign STORE_DATA_PORT_LSQ_dist_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 79:31:@14698.4]
  assign STORE_ADDR_PORT_LSQ_dist_clock = clock; // @[:@14703.4]
  assign STORE_ADDR_PORT_LSQ_dist_reset = reset; // @[:@14704.4]
  assign STORE_ADDR_PORT_LSQ_dist_io_dataFromPrev_valid = io_wrAddrPorts_0_valid; // @[LSQBRAM.scala 82:34:@14710.4]
  assign STORE_ADDR_PORT_LSQ_dist_io_dataFromPrev_bits = io_wrAddrPorts_0_bits; // @[LSQBRAM.scala 82:34:@14709.4]
  assign STORE_ADDR_PORT_LSQ_dist_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 82:34:@14708.4]
endmodule
