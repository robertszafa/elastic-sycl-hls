module STORE_QUEUE_LSQ_A( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_bbStart, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_0, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_1, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_2, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_3, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_4, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_5, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_6, // @[:@6.4]
  input  [2:0]  io_bbStoreOffsets_7, // @[:@6.4]
  input         io_bbStorePorts_1, // @[:@6.4]
  input  [1:0]  io_bbNumStores, // @[:@6.4]
  output [2:0]  io_storeTail, // @[:@6.4]
  output [2:0]  io_storeHead, // @[:@6.4]
  output        io_storeEmpty, // @[:@6.4]
  input  [2:0]  io_loadTail, // @[:@6.4]
  input  [2:0]  io_loadHead, // @[:@6.4]
  input         io_loadEmpty, // @[:@6.4]
  input         io_loadAddressDone_0, // @[:@6.4]
  input         io_loadAddressDone_1, // @[:@6.4]
  input         io_loadAddressDone_2, // @[:@6.4]
  input         io_loadAddressDone_3, // @[:@6.4]
  input         io_loadAddressDone_4, // @[:@6.4]
  input         io_loadAddressDone_5, // @[:@6.4]
  input         io_loadAddressDone_6, // @[:@6.4]
  input         io_loadAddressDone_7, // @[:@6.4]
  input         io_loadDataDone_0, // @[:@6.4]
  input         io_loadDataDone_1, // @[:@6.4]
  input         io_loadDataDone_2, // @[:@6.4]
  input         io_loadDataDone_3, // @[:@6.4]
  input         io_loadDataDone_4, // @[:@6.4]
  input         io_loadDataDone_5, // @[:@6.4]
  input         io_loadDataDone_6, // @[:@6.4]
  input         io_loadDataDone_7, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_0, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_1, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_2, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_3, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_4, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_5, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_6, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_7, // @[:@6.4]
  output        io_storeAddrDone_0, // @[:@6.4]
  output        io_storeAddrDone_1, // @[:@6.4]
  output        io_storeAddrDone_2, // @[:@6.4]
  output        io_storeAddrDone_3, // @[:@6.4]
  output        io_storeAddrDone_4, // @[:@6.4]
  output        io_storeAddrDone_5, // @[:@6.4]
  output        io_storeAddrDone_6, // @[:@6.4]
  output        io_storeAddrDone_7, // @[:@6.4]
  output        io_storeDataDone_0, // @[:@6.4]
  output        io_storeDataDone_1, // @[:@6.4]
  output        io_storeDataDone_2, // @[:@6.4]
  output        io_storeDataDone_3, // @[:@6.4]
  output        io_storeDataDone_4, // @[:@6.4]
  output        io_storeDataDone_5, // @[:@6.4]
  output        io_storeDataDone_6, // @[:@6.4]
  output        io_storeDataDone_7, // @[:@6.4]
  output [31:0] io_storeAddrQueue_0, // @[:@6.4]
  output [31:0] io_storeAddrQueue_1, // @[:@6.4]
  output [31:0] io_storeAddrQueue_2, // @[:@6.4]
  output [31:0] io_storeAddrQueue_3, // @[:@6.4]
  output [31:0] io_storeAddrQueue_4, // @[:@6.4]
  output [31:0] io_storeAddrQueue_5, // @[:@6.4]
  output [31:0] io_storeAddrQueue_6, // @[:@6.4]
  output [31:0] io_storeAddrQueue_7, // @[:@6.4]
  output [31:0] io_storeDataQueue_0, // @[:@6.4]
  output [31:0] io_storeDataQueue_1, // @[:@6.4]
  output [31:0] io_storeDataQueue_2, // @[:@6.4]
  output [31:0] io_storeDataQueue_3, // @[:@6.4]
  output [31:0] io_storeDataQueue_4, // @[:@6.4]
  output [31:0] io_storeDataQueue_5, // @[:@6.4]
  output [31:0] io_storeDataQueue_6, // @[:@6.4]
  output [31:0] io_storeDataQueue_7, // @[:@6.4]
  input         io_storeDataEnable_0, // @[:@6.4]
  input         io_storeDataEnable_1, // @[:@6.4]
  input  [31:0] io_dataFromStorePorts_0, // @[:@6.4]
  input  [31:0] io_dataFromStorePorts_1, // @[:@6.4]
  input         io_storeAddrEnable_0, // @[:@6.4]
  input         io_storeAddrEnable_1, // @[:@6.4]
  input  [31:0] io_addressFromStorePorts_0, // @[:@6.4]
  input  [31:0] io_addressFromStorePorts_1, // @[:@6.4]
  output [31:0] io_storeAddrToMem, // @[:@6.4]
  output [31:0] io_storeDataToMem, // @[:@6.4]
  output        io_storeEnableToMem, // @[:@6.4]
  input         io_memIsReadyForStores // @[:@6.4]
);
  reg [2:0] head; // @[StoreQueue.scala 50:21:@8.4]
  reg [31:0] _RAND_0;
  reg [2:0] tail; // @[StoreQueue.scala 51:21:@9.4]
  reg [31:0] _RAND_1;
  reg [2:0] offsetQ_0; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_2;
  reg [2:0] offsetQ_1; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_3;
  reg [2:0] offsetQ_2; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_4;
  reg [2:0] offsetQ_3; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_5;
  reg [2:0] offsetQ_4; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_6;
  reg [2:0] offsetQ_5; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_7;
  reg [2:0] offsetQ_6; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_8;
  reg [2:0] offsetQ_7; // @[StoreQueue.scala 53:24:@19.4]
  reg [31:0] _RAND_9;
  reg  portQ_0; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_10;
  reg  portQ_1; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_11;
  reg  portQ_2; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_12;
  reg  portQ_3; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_13;
  reg  portQ_4; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_14;
  reg  portQ_5; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_15;
  reg  portQ_6; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_16;
  reg  portQ_7; // @[StoreQueue.scala 54:22:@29.4]
  reg [31:0] _RAND_17;
  reg [31:0] addrQ_0; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_18;
  reg [31:0] addrQ_1; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_19;
  reg [31:0] addrQ_2; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_20;
  reg [31:0] addrQ_3; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_21;
  reg [31:0] addrQ_4; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_22;
  reg [31:0] addrQ_5; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_23;
  reg [31:0] addrQ_6; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_24;
  reg [31:0] addrQ_7; // @[StoreQueue.scala 55:22:@39.4]
  reg [31:0] _RAND_25;
  reg [31:0] dataQ_0; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_26;
  reg [31:0] dataQ_1; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_27;
  reg [31:0] dataQ_2; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_28;
  reg [31:0] dataQ_3; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_29;
  reg [31:0] dataQ_4; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_30;
  reg [31:0] dataQ_5; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_31;
  reg [31:0] dataQ_6; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_32;
  reg [31:0] dataQ_7; // @[StoreQueue.scala 56:22:@49.4]
  reg [31:0] _RAND_33;
  reg  addrKnown_0; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_34;
  reg  addrKnown_1; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_35;
  reg  addrKnown_2; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_36;
  reg  addrKnown_3; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_37;
  reg  addrKnown_4; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_38;
  reg  addrKnown_5; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_39;
  reg  addrKnown_6; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_40;
  reg  addrKnown_7; // @[StoreQueue.scala 57:26:@59.4]
  reg [31:0] _RAND_41;
  reg  dataKnown_0; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_42;
  reg  dataKnown_1; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_43;
  reg  dataKnown_2; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_44;
  reg  dataKnown_3; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_45;
  reg  dataKnown_4; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_46;
  reg  dataKnown_5; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_47;
  reg  dataKnown_6; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_48;
  reg  dataKnown_7; // @[StoreQueue.scala 58:26:@69.4]
  reg [31:0] _RAND_49;
  reg  allocatedEntries_0; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_50;
  reg  allocatedEntries_1; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_51;
  reg  allocatedEntries_2; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_52;
  reg  allocatedEntries_3; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_53;
  reg  allocatedEntries_4; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_54;
  reg  allocatedEntries_5; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_55;
  reg  allocatedEntries_6; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_56;
  reg  allocatedEntries_7; // @[StoreQueue.scala 59:33:@79.4]
  reg [31:0] _RAND_57;
  reg  storeCompleted_0; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_58;
  reg  storeCompleted_1; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_59;
  reg  storeCompleted_2; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_60;
  reg  storeCompleted_3; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_61;
  reg  storeCompleted_4; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_62;
  reg  storeCompleted_5; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_63;
  reg  storeCompleted_6; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_64;
  reg  storeCompleted_7; // @[StoreQueue.scala 60:31:@89.4]
  reg [31:0] _RAND_65;
  reg  checkBits_0; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_66;
  reg  checkBits_1; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_67;
  reg  checkBits_2; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_68;
  reg  checkBits_3; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_69;
  reg  checkBits_4; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_70;
  reg  checkBits_5; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_71;
  reg  checkBits_6; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_72;
  reg  checkBits_7; // @[StoreQueue.scala 61:26:@99.4]
  reg [31:0] _RAND_73;
  wire [4:0] _GEN_410; // @[util.scala 14:20:@101.4]
  wire [5:0] _T_956; // @[util.scala 14:20:@101.4]
  wire [5:0] _T_957; // @[util.scala 14:20:@102.4]
  wire [4:0] _T_958; // @[util.scala 14:20:@103.4]
  wire [4:0] _GEN_0; // @[util.scala 14:25:@104.4]
  wire [3:0] _T_959; // @[util.scala 14:25:@104.4]
  wire [3:0] _GEN_411; // @[StoreQueue.scala 70:46:@105.4]
  wire  _T_960; // @[StoreQueue.scala 70:46:@105.4]
  wire  initBits_0; // @[StoreQueue.scala 70:64:@106.4]
  wire [5:0] _T_965; // @[util.scala 14:20:@108.4]
  wire [5:0] _T_966; // @[util.scala 14:20:@109.4]
  wire [4:0] _T_967; // @[util.scala 14:20:@110.4]
  wire [4:0] _GEN_8; // @[util.scala 14:25:@111.4]
  wire [3:0] _T_968; // @[util.scala 14:25:@111.4]
  wire  _T_969; // @[StoreQueue.scala 70:46:@112.4]
  wire  initBits_1; // @[StoreQueue.scala 70:64:@113.4]
  wire [5:0] _T_974; // @[util.scala 14:20:@115.4]
  wire [5:0] _T_975; // @[util.scala 14:20:@116.4]
  wire [4:0] _T_976; // @[util.scala 14:20:@117.4]
  wire [4:0] _GEN_18; // @[util.scala 14:25:@118.4]
  wire [3:0] _T_977; // @[util.scala 14:25:@118.4]
  wire  _T_978; // @[StoreQueue.scala 70:46:@119.4]
  wire  initBits_2; // @[StoreQueue.scala 70:64:@120.4]
  wire [5:0] _T_983; // @[util.scala 14:20:@122.4]
  wire [5:0] _T_984; // @[util.scala 14:20:@123.4]
  wire [4:0] _T_985; // @[util.scala 14:20:@124.4]
  wire [4:0] _GEN_26; // @[util.scala 14:25:@125.4]
  wire [3:0] _T_986; // @[util.scala 14:25:@125.4]
  wire  _T_987; // @[StoreQueue.scala 70:46:@126.4]
  wire  initBits_3; // @[StoreQueue.scala 70:64:@127.4]
  wire [5:0] _T_992; // @[util.scala 14:20:@129.4]
  wire [5:0] _T_993; // @[util.scala 14:20:@130.4]
  wire [4:0] _T_994; // @[util.scala 14:20:@131.4]
  wire [4:0] _GEN_36; // @[util.scala 14:25:@132.4]
  wire [3:0] _T_995; // @[util.scala 14:25:@132.4]
  wire  _T_996; // @[StoreQueue.scala 70:46:@133.4]
  wire  initBits_4; // @[StoreQueue.scala 70:64:@134.4]
  wire [5:0] _T_1001; // @[util.scala 14:20:@136.4]
  wire [5:0] _T_1002; // @[util.scala 14:20:@137.4]
  wire [4:0] _T_1003; // @[util.scala 14:20:@138.4]
  wire [4:0] _GEN_44; // @[util.scala 14:25:@139.4]
  wire [3:0] _T_1004; // @[util.scala 14:25:@139.4]
  wire  _T_1005; // @[StoreQueue.scala 70:46:@140.4]
  wire  initBits_5; // @[StoreQueue.scala 70:64:@141.4]
  wire [5:0] _T_1010; // @[util.scala 14:20:@143.4]
  wire [5:0] _T_1011; // @[util.scala 14:20:@144.4]
  wire [4:0] _T_1012; // @[util.scala 14:20:@145.4]
  wire [4:0] _GEN_54; // @[util.scala 14:25:@146.4]
  wire [3:0] _T_1013; // @[util.scala 14:25:@146.4]
  wire  _T_1014; // @[StoreQueue.scala 70:46:@147.4]
  wire  initBits_6; // @[StoreQueue.scala 70:64:@148.4]
  wire [5:0] _T_1019; // @[util.scala 14:20:@150.4]
  wire [5:0] _T_1020; // @[util.scala 14:20:@151.4]
  wire [4:0] _T_1021; // @[util.scala 14:20:@152.4]
  wire [4:0] _GEN_62; // @[util.scala 14:25:@153.4]
  wire [3:0] _T_1022; // @[util.scala 14:25:@153.4]
  wire  _T_1023; // @[StoreQueue.scala 70:46:@154.4]
  wire  initBits_7; // @[StoreQueue.scala 70:64:@155.4]
  wire  _T_1038; // @[StoreQueue.scala 72:78:@165.4]
  wire  _T_1039; // @[StoreQueue.scala 72:78:@166.4]
  wire  _T_1040; // @[StoreQueue.scala 72:78:@167.4]
  wire  _T_1041; // @[StoreQueue.scala 72:78:@168.4]
  wire  _T_1042; // @[StoreQueue.scala 72:78:@169.4]
  wire  _T_1043; // @[StoreQueue.scala 72:78:@170.4]
  wire  _T_1044; // @[StoreQueue.scala 72:78:@171.4]
  wire  _T_1045; // @[StoreQueue.scala 72:78:@172.4]
  wire [2:0] _T_1068; // @[:@196.6]
  wire [2:0] _GEN_1; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_2; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_3; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_4; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_5; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_6; // @[StoreQueue.scala 76:20:@197.6]
  wire [2:0] _GEN_7; // @[StoreQueue.scala 76:20:@197.6]
  wire  _GEN_9; // @[StoreQueue.scala 77:18:@204.6]
  wire  _GEN_10; // @[StoreQueue.scala 77:18:@204.6]
  wire  _GEN_11; // @[StoreQueue.scala 77:18:@204.6]
  wire  _GEN_12; // @[StoreQueue.scala 77:18:@204.6]
  wire  _GEN_13; // @[StoreQueue.scala 77:18:@204.6]
  wire  _GEN_14; // @[StoreQueue.scala 77:18:@204.6]
  wire  _GEN_15; // @[StoreQueue.scala 77:18:@204.6]
  wire [2:0] _GEN_16; // @[StoreQueue.scala 75:25:@190.4]
  wire  _GEN_17; // @[StoreQueue.scala 75:25:@190.4]
  wire [2:0] _T_1086; // @[:@212.6]
  wire [2:0] _GEN_19; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_20; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_21; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_22; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_23; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_24; // @[StoreQueue.scala 76:20:@213.6]
  wire [2:0] _GEN_25; // @[StoreQueue.scala 76:20:@213.6]
  wire  _GEN_27; // @[StoreQueue.scala 77:18:@220.6]
  wire  _GEN_28; // @[StoreQueue.scala 77:18:@220.6]
  wire  _GEN_29; // @[StoreQueue.scala 77:18:@220.6]
  wire  _GEN_30; // @[StoreQueue.scala 77:18:@220.6]
  wire  _GEN_31; // @[StoreQueue.scala 77:18:@220.6]
  wire  _GEN_32; // @[StoreQueue.scala 77:18:@220.6]
  wire  _GEN_33; // @[StoreQueue.scala 77:18:@220.6]
  wire [2:0] _GEN_34; // @[StoreQueue.scala 75:25:@206.4]
  wire  _GEN_35; // @[StoreQueue.scala 75:25:@206.4]
  wire [2:0] _T_1104; // @[:@228.6]
  wire [2:0] _GEN_37; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_38; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_39; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_40; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_41; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_42; // @[StoreQueue.scala 76:20:@229.6]
  wire [2:0] _GEN_43; // @[StoreQueue.scala 76:20:@229.6]
  wire  _GEN_45; // @[StoreQueue.scala 77:18:@236.6]
  wire  _GEN_46; // @[StoreQueue.scala 77:18:@236.6]
  wire  _GEN_47; // @[StoreQueue.scala 77:18:@236.6]
  wire  _GEN_48; // @[StoreQueue.scala 77:18:@236.6]
  wire  _GEN_49; // @[StoreQueue.scala 77:18:@236.6]
  wire  _GEN_50; // @[StoreQueue.scala 77:18:@236.6]
  wire  _GEN_51; // @[StoreQueue.scala 77:18:@236.6]
  wire [2:0] _GEN_52; // @[StoreQueue.scala 75:25:@222.4]
  wire  _GEN_53; // @[StoreQueue.scala 75:25:@222.4]
  wire [2:0] _T_1122; // @[:@244.6]
  wire [2:0] _GEN_55; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_56; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_57; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_58; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_59; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_60; // @[StoreQueue.scala 76:20:@245.6]
  wire [2:0] _GEN_61; // @[StoreQueue.scala 76:20:@245.6]
  wire  _GEN_63; // @[StoreQueue.scala 77:18:@252.6]
  wire  _GEN_64; // @[StoreQueue.scala 77:18:@252.6]
  wire  _GEN_65; // @[StoreQueue.scala 77:18:@252.6]
  wire  _GEN_66; // @[StoreQueue.scala 77:18:@252.6]
  wire  _GEN_67; // @[StoreQueue.scala 77:18:@252.6]
  wire  _GEN_68; // @[StoreQueue.scala 77:18:@252.6]
  wire  _GEN_69; // @[StoreQueue.scala 77:18:@252.6]
  wire [2:0] _GEN_70; // @[StoreQueue.scala 75:25:@238.4]
  wire  _GEN_71; // @[StoreQueue.scala 75:25:@238.4]
  wire [2:0] _T_1140; // @[:@260.6]
  wire [2:0] _GEN_73; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_74; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_75; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_76; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_77; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_78; // @[StoreQueue.scala 76:20:@261.6]
  wire [2:0] _GEN_79; // @[StoreQueue.scala 76:20:@261.6]
  wire  _GEN_81; // @[StoreQueue.scala 77:18:@268.6]
  wire  _GEN_82; // @[StoreQueue.scala 77:18:@268.6]
  wire  _GEN_83; // @[StoreQueue.scala 77:18:@268.6]
  wire  _GEN_84; // @[StoreQueue.scala 77:18:@268.6]
  wire  _GEN_85; // @[StoreQueue.scala 77:18:@268.6]
  wire  _GEN_86; // @[StoreQueue.scala 77:18:@268.6]
  wire  _GEN_87; // @[StoreQueue.scala 77:18:@268.6]
  wire [2:0] _GEN_88; // @[StoreQueue.scala 75:25:@254.4]
  wire  _GEN_89; // @[StoreQueue.scala 75:25:@254.4]
  wire [2:0] _T_1158; // @[:@276.6]
  wire [2:0] _GEN_91; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_92; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_93; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_94; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_95; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_96; // @[StoreQueue.scala 76:20:@277.6]
  wire [2:0] _GEN_97; // @[StoreQueue.scala 76:20:@277.6]
  wire  _GEN_99; // @[StoreQueue.scala 77:18:@284.6]
  wire  _GEN_100; // @[StoreQueue.scala 77:18:@284.6]
  wire  _GEN_101; // @[StoreQueue.scala 77:18:@284.6]
  wire  _GEN_102; // @[StoreQueue.scala 77:18:@284.6]
  wire  _GEN_103; // @[StoreQueue.scala 77:18:@284.6]
  wire  _GEN_104; // @[StoreQueue.scala 77:18:@284.6]
  wire  _GEN_105; // @[StoreQueue.scala 77:18:@284.6]
  wire [2:0] _GEN_106; // @[StoreQueue.scala 75:25:@270.4]
  wire  _GEN_107; // @[StoreQueue.scala 75:25:@270.4]
  wire [2:0] _T_1176; // @[:@292.6]
  wire [2:0] _GEN_109; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_110; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_111; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_112; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_113; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_114; // @[StoreQueue.scala 76:20:@293.6]
  wire [2:0] _GEN_115; // @[StoreQueue.scala 76:20:@293.6]
  wire  _GEN_117; // @[StoreQueue.scala 77:18:@300.6]
  wire  _GEN_118; // @[StoreQueue.scala 77:18:@300.6]
  wire  _GEN_119; // @[StoreQueue.scala 77:18:@300.6]
  wire  _GEN_120; // @[StoreQueue.scala 77:18:@300.6]
  wire  _GEN_121; // @[StoreQueue.scala 77:18:@300.6]
  wire  _GEN_122; // @[StoreQueue.scala 77:18:@300.6]
  wire  _GEN_123; // @[StoreQueue.scala 77:18:@300.6]
  wire [2:0] _GEN_124; // @[StoreQueue.scala 75:25:@286.4]
  wire  _GEN_125; // @[StoreQueue.scala 75:25:@286.4]
  wire [2:0] _T_1194; // @[:@308.6]
  wire [2:0] _GEN_127; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_128; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_129; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_130; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_131; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_132; // @[StoreQueue.scala 76:20:@309.6]
  wire [2:0] _GEN_133; // @[StoreQueue.scala 76:20:@309.6]
  wire  _GEN_135; // @[StoreQueue.scala 77:18:@316.6]
  wire  _GEN_136; // @[StoreQueue.scala 77:18:@316.6]
  wire  _GEN_137; // @[StoreQueue.scala 77:18:@316.6]
  wire  _GEN_138; // @[StoreQueue.scala 77:18:@316.6]
  wire  _GEN_139; // @[StoreQueue.scala 77:18:@316.6]
  wire  _GEN_140; // @[StoreQueue.scala 77:18:@316.6]
  wire  _GEN_141; // @[StoreQueue.scala 77:18:@316.6]
  wire [2:0] _GEN_142; // @[StoreQueue.scala 75:25:@302.4]
  wire  _GEN_143; // @[StoreQueue.scala 75:25:@302.4]
  reg [2:0] previousLoadHead; // @[StoreQueue.scala 92:33:@318.4]
  reg [31:0] _RAND_74;
  wire [3:0] _T_1216; // @[util.scala 10:8:@327.6]
  wire [3:0] _GEN_72; // @[util.scala 10:14:@328.6]
  wire [3:0] _T_1217; // @[util.scala 10:14:@328.6]
  wire [3:0] _GEN_443; // @[StoreQueue.scala 96:56:@329.6]
  wire  _T_1218; // @[StoreQueue.scala 96:56:@329.6]
  wire  _T_1219; // @[StoreQueue.scala 95:50:@330.6]
  wire  _T_1221; // @[StoreQueue.scala 95:35:@331.6]
  wire  _T_1223; // @[StoreQueue.scala 100:35:@339.8]
  wire  _T_1224; // @[StoreQueue.scala 100:87:@340.8]
  wire  _T_1225; // @[StoreQueue.scala 100:61:@341.8]
  wire  _T_1227; // @[StoreQueue.scala 102:35:@346.10]
  wire  _T_1228; // @[StoreQueue.scala 103:23:@347.10]
  wire  _T_1229; // @[StoreQueue.scala 103:75:@348.10]
  wire  _T_1230; // @[StoreQueue.scala 103:49:@349.10]
  wire  _T_1232; // @[StoreQueue.scala 103:9:@350.10]
  wire  _T_1233; // @[StoreQueue.scala 102:49:@351.10]
  wire  _GEN_152; // @[StoreQueue.scala 103:96:@352.10]
  wire  _GEN_153; // @[StoreQueue.scala 100:102:@342.8]
  wire  _GEN_154; // @[StoreQueue.scala 98:26:@335.6]
  wire  _GEN_155; // @[StoreQueue.scala 94:35:@320.4]
  wire [3:0] _T_1246; // @[util.scala 10:8:@363.6]
  wire [3:0] _GEN_80; // @[util.scala 10:14:@364.6]
  wire [3:0] _T_1247; // @[util.scala 10:14:@364.6]
  wire  _T_1248; // @[StoreQueue.scala 96:56:@365.6]
  wire  _T_1249; // @[StoreQueue.scala 95:50:@366.6]
  wire  _T_1251; // @[StoreQueue.scala 95:35:@367.6]
  wire  _T_1253; // @[StoreQueue.scala 100:35:@375.8]
  wire  _T_1254; // @[StoreQueue.scala 100:87:@376.8]
  wire  _T_1255; // @[StoreQueue.scala 100:61:@377.8]
  wire  _T_1258; // @[StoreQueue.scala 103:23:@383.10]
  wire  _T_1259; // @[StoreQueue.scala 103:75:@384.10]
  wire  _T_1260; // @[StoreQueue.scala 103:49:@385.10]
  wire  _T_1262; // @[StoreQueue.scala 103:9:@386.10]
  wire  _T_1263; // @[StoreQueue.scala 102:49:@387.10]
  wire  _GEN_164; // @[StoreQueue.scala 103:96:@388.10]
  wire  _GEN_165; // @[StoreQueue.scala 100:102:@378.8]
  wire  _GEN_166; // @[StoreQueue.scala 98:26:@371.6]
  wire  _GEN_167; // @[StoreQueue.scala 94:35:@356.4]
  wire [3:0] _T_1276; // @[util.scala 10:8:@399.6]
  wire [3:0] _GEN_90; // @[util.scala 10:14:@400.6]
  wire [3:0] _T_1277; // @[util.scala 10:14:@400.6]
  wire  _T_1278; // @[StoreQueue.scala 96:56:@401.6]
  wire  _T_1279; // @[StoreQueue.scala 95:50:@402.6]
  wire  _T_1281; // @[StoreQueue.scala 95:35:@403.6]
  wire  _T_1283; // @[StoreQueue.scala 100:35:@411.8]
  wire  _T_1284; // @[StoreQueue.scala 100:87:@412.8]
  wire  _T_1285; // @[StoreQueue.scala 100:61:@413.8]
  wire  _T_1288; // @[StoreQueue.scala 103:23:@419.10]
  wire  _T_1289; // @[StoreQueue.scala 103:75:@420.10]
  wire  _T_1290; // @[StoreQueue.scala 103:49:@421.10]
  wire  _T_1292; // @[StoreQueue.scala 103:9:@422.10]
  wire  _T_1293; // @[StoreQueue.scala 102:49:@423.10]
  wire  _GEN_176; // @[StoreQueue.scala 103:96:@424.10]
  wire  _GEN_177; // @[StoreQueue.scala 100:102:@414.8]
  wire  _GEN_178; // @[StoreQueue.scala 98:26:@407.6]
  wire  _GEN_179; // @[StoreQueue.scala 94:35:@392.4]
  wire [3:0] _T_1306; // @[util.scala 10:8:@435.6]
  wire [3:0] _GEN_98; // @[util.scala 10:14:@436.6]
  wire [3:0] _T_1307; // @[util.scala 10:14:@436.6]
  wire  _T_1308; // @[StoreQueue.scala 96:56:@437.6]
  wire  _T_1309; // @[StoreQueue.scala 95:50:@438.6]
  wire  _T_1311; // @[StoreQueue.scala 95:35:@439.6]
  wire  _T_1313; // @[StoreQueue.scala 100:35:@447.8]
  wire  _T_1314; // @[StoreQueue.scala 100:87:@448.8]
  wire  _T_1315; // @[StoreQueue.scala 100:61:@449.8]
  wire  _T_1318; // @[StoreQueue.scala 103:23:@455.10]
  wire  _T_1319; // @[StoreQueue.scala 103:75:@456.10]
  wire  _T_1320; // @[StoreQueue.scala 103:49:@457.10]
  wire  _T_1322; // @[StoreQueue.scala 103:9:@458.10]
  wire  _T_1323; // @[StoreQueue.scala 102:49:@459.10]
  wire  _GEN_188; // @[StoreQueue.scala 103:96:@460.10]
  wire  _GEN_189; // @[StoreQueue.scala 100:102:@450.8]
  wire  _GEN_190; // @[StoreQueue.scala 98:26:@443.6]
  wire  _GEN_191; // @[StoreQueue.scala 94:35:@428.4]
  wire [3:0] _T_1336; // @[util.scala 10:8:@471.6]
  wire [3:0] _GEN_108; // @[util.scala 10:14:@472.6]
  wire [3:0] _T_1337; // @[util.scala 10:14:@472.6]
  wire  _T_1338; // @[StoreQueue.scala 96:56:@473.6]
  wire  _T_1339; // @[StoreQueue.scala 95:50:@474.6]
  wire  _T_1341; // @[StoreQueue.scala 95:35:@475.6]
  wire  _T_1343; // @[StoreQueue.scala 100:35:@483.8]
  wire  _T_1344; // @[StoreQueue.scala 100:87:@484.8]
  wire  _T_1345; // @[StoreQueue.scala 100:61:@485.8]
  wire  _T_1348; // @[StoreQueue.scala 103:23:@491.10]
  wire  _T_1349; // @[StoreQueue.scala 103:75:@492.10]
  wire  _T_1350; // @[StoreQueue.scala 103:49:@493.10]
  wire  _T_1352; // @[StoreQueue.scala 103:9:@494.10]
  wire  _T_1353; // @[StoreQueue.scala 102:49:@495.10]
  wire  _GEN_200; // @[StoreQueue.scala 103:96:@496.10]
  wire  _GEN_201; // @[StoreQueue.scala 100:102:@486.8]
  wire  _GEN_202; // @[StoreQueue.scala 98:26:@479.6]
  wire  _GEN_203; // @[StoreQueue.scala 94:35:@464.4]
  wire [3:0] _T_1366; // @[util.scala 10:8:@507.6]
  wire [3:0] _GEN_116; // @[util.scala 10:14:@508.6]
  wire [3:0] _T_1367; // @[util.scala 10:14:@508.6]
  wire  _T_1368; // @[StoreQueue.scala 96:56:@509.6]
  wire  _T_1369; // @[StoreQueue.scala 95:50:@510.6]
  wire  _T_1371; // @[StoreQueue.scala 95:35:@511.6]
  wire  _T_1373; // @[StoreQueue.scala 100:35:@519.8]
  wire  _T_1374; // @[StoreQueue.scala 100:87:@520.8]
  wire  _T_1375; // @[StoreQueue.scala 100:61:@521.8]
  wire  _T_1378; // @[StoreQueue.scala 103:23:@527.10]
  wire  _T_1379; // @[StoreQueue.scala 103:75:@528.10]
  wire  _T_1380; // @[StoreQueue.scala 103:49:@529.10]
  wire  _T_1382; // @[StoreQueue.scala 103:9:@530.10]
  wire  _T_1383; // @[StoreQueue.scala 102:49:@531.10]
  wire  _GEN_212; // @[StoreQueue.scala 103:96:@532.10]
  wire  _GEN_213; // @[StoreQueue.scala 100:102:@522.8]
  wire  _GEN_214; // @[StoreQueue.scala 98:26:@515.6]
  wire  _GEN_215; // @[StoreQueue.scala 94:35:@500.4]
  wire [3:0] _T_1396; // @[util.scala 10:8:@543.6]
  wire [3:0] _GEN_126; // @[util.scala 10:14:@544.6]
  wire [3:0] _T_1397; // @[util.scala 10:14:@544.6]
  wire  _T_1398; // @[StoreQueue.scala 96:56:@545.6]
  wire  _T_1399; // @[StoreQueue.scala 95:50:@546.6]
  wire  _T_1401; // @[StoreQueue.scala 95:35:@547.6]
  wire  _T_1403; // @[StoreQueue.scala 100:35:@555.8]
  wire  _T_1404; // @[StoreQueue.scala 100:87:@556.8]
  wire  _T_1405; // @[StoreQueue.scala 100:61:@557.8]
  wire  _T_1408; // @[StoreQueue.scala 103:23:@563.10]
  wire  _T_1409; // @[StoreQueue.scala 103:75:@564.10]
  wire  _T_1410; // @[StoreQueue.scala 103:49:@565.10]
  wire  _T_1412; // @[StoreQueue.scala 103:9:@566.10]
  wire  _T_1413; // @[StoreQueue.scala 102:49:@567.10]
  wire  _GEN_224; // @[StoreQueue.scala 103:96:@568.10]
  wire  _GEN_225; // @[StoreQueue.scala 100:102:@558.8]
  wire  _GEN_226; // @[StoreQueue.scala 98:26:@551.6]
  wire  _GEN_227; // @[StoreQueue.scala 94:35:@536.4]
  wire [3:0] _T_1426; // @[util.scala 10:8:@579.6]
  wire [3:0] _GEN_134; // @[util.scala 10:14:@580.6]
  wire [3:0] _T_1427; // @[util.scala 10:14:@580.6]
  wire  _T_1428; // @[StoreQueue.scala 96:56:@581.6]
  wire  _T_1429; // @[StoreQueue.scala 95:50:@582.6]
  wire  _T_1431; // @[StoreQueue.scala 95:35:@583.6]
  wire  _T_1433; // @[StoreQueue.scala 100:35:@591.8]
  wire  _T_1434; // @[StoreQueue.scala 100:87:@592.8]
  wire  _T_1435; // @[StoreQueue.scala 100:61:@593.8]
  wire  _T_1438; // @[StoreQueue.scala 103:23:@599.10]
  wire  _T_1439; // @[StoreQueue.scala 103:75:@600.10]
  wire  _T_1440; // @[StoreQueue.scala 103:49:@601.10]
  wire  _T_1442; // @[StoreQueue.scala 103:9:@602.10]
  wire  _T_1443; // @[StoreQueue.scala 102:49:@603.10]
  wire  _GEN_236; // @[StoreQueue.scala 103:96:@604.10]
  wire  _GEN_237; // @[StoreQueue.scala 100:102:@594.8]
  wire  _GEN_238; // @[StoreQueue.scala 98:26:@587.6]
  wire  _GEN_239; // @[StoreQueue.scala 94:35:@572.4]
  wire  _T_1445; // @[StoreQueue.scala 119:103:@608.4]
  wire  _T_1447; // @[StoreQueue.scala 120:17:@609.4]
  wire  _T_1449; // @[StoreQueue.scala 120:35:@610.4]
  wire  _T_1450; // @[StoreQueue.scala 120:26:@611.4]
  wire  _T_1452; // @[StoreQueue.scala 120:50:@612.4]
  wire  _T_1454; // @[StoreQueue.scala 120:81:@613.4]
  wire  _T_1456; // @[StoreQueue.scala 120:99:@614.4]
  wire  _T_1457; // @[StoreQueue.scala 120:90:@615.4]
  wire  _T_1459; // @[StoreQueue.scala 120:67:@616.4]
  wire  _T_1460; // @[StoreQueue.scala 120:64:@617.4]
  wire  validEntriesInLoadQ_0; // @[StoreQueue.scala 119:90:@618.4]
  wire  _T_1464; // @[StoreQueue.scala 120:17:@620.4]
  wire  _T_1466; // @[StoreQueue.scala 120:35:@621.4]
  wire  _T_1467; // @[StoreQueue.scala 120:26:@622.4]
  wire  _T_1471; // @[StoreQueue.scala 120:81:@624.4]
  wire  _T_1473; // @[StoreQueue.scala 120:99:@625.4]
  wire  _T_1474; // @[StoreQueue.scala 120:90:@626.4]
  wire  _T_1476; // @[StoreQueue.scala 120:67:@627.4]
  wire  _T_1477; // @[StoreQueue.scala 120:64:@628.4]
  wire  validEntriesInLoadQ_1; // @[StoreQueue.scala 119:90:@629.4]
  wire  _T_1481; // @[StoreQueue.scala 120:17:@631.4]
  wire  _T_1483; // @[StoreQueue.scala 120:35:@632.4]
  wire  _T_1484; // @[StoreQueue.scala 120:26:@633.4]
  wire  _T_1488; // @[StoreQueue.scala 120:81:@635.4]
  wire  _T_1490; // @[StoreQueue.scala 120:99:@636.4]
  wire  _T_1491; // @[StoreQueue.scala 120:90:@637.4]
  wire  _T_1493; // @[StoreQueue.scala 120:67:@638.4]
  wire  _T_1494; // @[StoreQueue.scala 120:64:@639.4]
  wire  validEntriesInLoadQ_2; // @[StoreQueue.scala 119:90:@640.4]
  wire  _T_1498; // @[StoreQueue.scala 120:17:@642.4]
  wire  _T_1500; // @[StoreQueue.scala 120:35:@643.4]
  wire  _T_1501; // @[StoreQueue.scala 120:26:@644.4]
  wire  _T_1505; // @[StoreQueue.scala 120:81:@646.4]
  wire  _T_1507; // @[StoreQueue.scala 120:99:@647.4]
  wire  _T_1508; // @[StoreQueue.scala 120:90:@648.4]
  wire  _T_1510; // @[StoreQueue.scala 120:67:@649.4]
  wire  _T_1511; // @[StoreQueue.scala 120:64:@650.4]
  wire  validEntriesInLoadQ_3; // @[StoreQueue.scala 119:90:@651.4]
  wire  _T_1515; // @[StoreQueue.scala 120:17:@653.4]
  wire  _T_1517; // @[StoreQueue.scala 120:35:@654.4]
  wire  _T_1518; // @[StoreQueue.scala 120:26:@655.4]
  wire  _T_1522; // @[StoreQueue.scala 120:81:@657.4]
  wire  _T_1524; // @[StoreQueue.scala 120:99:@658.4]
  wire  _T_1525; // @[StoreQueue.scala 120:90:@659.4]
  wire  _T_1527; // @[StoreQueue.scala 120:67:@660.4]
  wire  _T_1528; // @[StoreQueue.scala 120:64:@661.4]
  wire  validEntriesInLoadQ_4; // @[StoreQueue.scala 119:90:@662.4]
  wire  _T_1532; // @[StoreQueue.scala 120:17:@664.4]
  wire  _T_1534; // @[StoreQueue.scala 120:35:@665.4]
  wire  _T_1535; // @[StoreQueue.scala 120:26:@666.4]
  wire  _T_1539; // @[StoreQueue.scala 120:81:@668.4]
  wire  _T_1541; // @[StoreQueue.scala 120:99:@669.4]
  wire  _T_1542; // @[StoreQueue.scala 120:90:@670.4]
  wire  _T_1544; // @[StoreQueue.scala 120:67:@671.4]
  wire  _T_1545; // @[StoreQueue.scala 120:64:@672.4]
  wire  validEntriesInLoadQ_5; // @[StoreQueue.scala 119:90:@673.4]
  wire  _T_1549; // @[StoreQueue.scala 120:17:@675.4]
  wire  _T_1551; // @[StoreQueue.scala 120:35:@676.4]
  wire  _T_1552; // @[StoreQueue.scala 120:26:@677.4]
  wire  _T_1556; // @[StoreQueue.scala 120:81:@679.4]
  wire  _T_1558; // @[StoreQueue.scala 120:99:@680.4]
  wire  _T_1559; // @[StoreQueue.scala 120:90:@681.4]
  wire  _T_1561; // @[StoreQueue.scala 120:67:@682.4]
  wire  _T_1562; // @[StoreQueue.scala 120:64:@683.4]
  wire  validEntriesInLoadQ_6; // @[StoreQueue.scala 119:90:@684.4]
  wire  validEntriesInLoadQ_7; // @[StoreQueue.scala 119:90:@695.4]
  wire [2:0] _GEN_241; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_242; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_243; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_244; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_245; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_246; // @[StoreQueue.scala 126:96:@705.4]
  wire [2:0] _GEN_247; // @[StoreQueue.scala 126:96:@705.4]
  wire  _T_1597; // @[StoreQueue.scala 126:96:@705.4]
  wire  loadsToCheck_0; // @[StoreQueue.scala 126:83:@713.4]
  wire  _T_1627; // @[StoreQueue.scala 127:37:@716.4]
  wire  _T_1628; // @[StoreQueue.scala 127:28:@717.4]
  wire  _T_1633; // @[StoreQueue.scala 127:71:@718.4]
  wire  _T_1636; // @[StoreQueue.scala 127:79:@720.4]
  wire  _T_1638; // @[StoreQueue.scala 127:55:@721.4]
  wire  loadsToCheck_1; // @[StoreQueue.scala 126:83:@722.4]
  wire  _T_1650; // @[StoreQueue.scala 127:37:@725.4]
  wire  _T_1651; // @[StoreQueue.scala 127:28:@726.4]
  wire  _T_1656; // @[StoreQueue.scala 127:71:@727.4]
  wire  _T_1659; // @[StoreQueue.scala 127:79:@729.4]
  wire  _T_1661; // @[StoreQueue.scala 127:55:@730.4]
  wire  loadsToCheck_2; // @[StoreQueue.scala 126:83:@731.4]
  wire  _T_1673; // @[StoreQueue.scala 127:37:@734.4]
  wire  _T_1674; // @[StoreQueue.scala 127:28:@735.4]
  wire  _T_1679; // @[StoreQueue.scala 127:71:@736.4]
  wire  _T_1682; // @[StoreQueue.scala 127:79:@738.4]
  wire  _T_1684; // @[StoreQueue.scala 127:55:@739.4]
  wire  loadsToCheck_3; // @[StoreQueue.scala 126:83:@740.4]
  wire  _T_1696; // @[StoreQueue.scala 127:37:@743.4]
  wire  _T_1697; // @[StoreQueue.scala 127:28:@744.4]
  wire  _T_1702; // @[StoreQueue.scala 127:71:@745.4]
  wire  _T_1705; // @[StoreQueue.scala 127:79:@747.4]
  wire  _T_1707; // @[StoreQueue.scala 127:55:@748.4]
  wire  loadsToCheck_4; // @[StoreQueue.scala 126:83:@749.4]
  wire  _T_1719; // @[StoreQueue.scala 127:37:@752.4]
  wire  _T_1720; // @[StoreQueue.scala 127:28:@753.4]
  wire  _T_1725; // @[StoreQueue.scala 127:71:@754.4]
  wire  _T_1728; // @[StoreQueue.scala 127:79:@756.4]
  wire  _T_1730; // @[StoreQueue.scala 127:55:@757.4]
  wire  loadsToCheck_5; // @[StoreQueue.scala 126:83:@758.4]
  wire  _T_1742; // @[StoreQueue.scala 127:37:@761.4]
  wire  _T_1743; // @[StoreQueue.scala 127:28:@762.4]
  wire  _T_1748; // @[StoreQueue.scala 127:71:@763.4]
  wire  _T_1751; // @[StoreQueue.scala 127:79:@765.4]
  wire  _T_1753; // @[StoreQueue.scala 127:55:@766.4]
  wire  loadsToCheck_6; // @[StoreQueue.scala 126:83:@767.4]
  wire  _T_1765; // @[StoreQueue.scala 127:37:@770.4]
  wire  loadsToCheck_7; // @[StoreQueue.scala 126:83:@776.4]
  wire  _T_1791; // @[StoreQueue.scala 133:16:@786.4]
  wire  _GEN_249; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_250; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_251; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_252; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_253; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_254; // @[StoreQueue.scala 133:24:@787.4]
  wire  _GEN_255; // @[StoreQueue.scala 133:24:@787.4]
  wire  entriesToCheck_0; // @[StoreQueue.scala 133:24:@787.4]
  wire  _T_1796; // @[StoreQueue.scala 133:16:@788.4]
  wire  entriesToCheck_1; // @[StoreQueue.scala 133:24:@789.4]
  wire  _T_1801; // @[StoreQueue.scala 133:16:@790.4]
  wire  entriesToCheck_2; // @[StoreQueue.scala 133:24:@791.4]
  wire  _T_1806; // @[StoreQueue.scala 133:16:@792.4]
  wire  entriesToCheck_3; // @[StoreQueue.scala 133:24:@793.4]
  wire  _T_1811; // @[StoreQueue.scala 133:16:@794.4]
  wire  entriesToCheck_4; // @[StoreQueue.scala 133:24:@795.4]
  wire  _T_1816; // @[StoreQueue.scala 133:16:@796.4]
  wire  entriesToCheck_5; // @[StoreQueue.scala 133:24:@797.4]
  wire  _T_1821; // @[StoreQueue.scala 133:16:@798.4]
  wire  entriesToCheck_6; // @[StoreQueue.scala 133:24:@799.4]
  wire  _T_1826; // @[StoreQueue.scala 133:16:@800.4]
  wire  entriesToCheck_7; // @[StoreQueue.scala 133:24:@801.4]
  wire  _T_1858; // @[StoreQueue.scala 140:34:@812.4]
  wire  _T_1859; // @[StoreQueue.scala 140:64:@813.4]
  wire [31:0] _GEN_257; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_258; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_259; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_260; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_261; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_262; // @[StoreQueue.scala 141:51:@814.4]
  wire [31:0] _GEN_263; // @[StoreQueue.scala 141:51:@814.4]
  wire  _T_1863; // @[StoreQueue.scala 141:51:@814.4]
  wire  _T_1864; // @[StoreQueue.scala 141:36:@815.4]
  wire  noConflicts_0; // @[StoreQueue.scala 140:95:@816.4]
  wire  _T_1867; // @[StoreQueue.scala 140:34:@818.4]
  wire  _T_1868; // @[StoreQueue.scala 140:64:@819.4]
  wire  _T_1872; // @[StoreQueue.scala 141:51:@820.4]
  wire  _T_1873; // @[StoreQueue.scala 141:36:@821.4]
  wire  noConflicts_1; // @[StoreQueue.scala 140:95:@822.4]
  wire  _T_1876; // @[StoreQueue.scala 140:34:@824.4]
  wire  _T_1877; // @[StoreQueue.scala 140:64:@825.4]
  wire  _T_1881; // @[StoreQueue.scala 141:51:@826.4]
  wire  _T_1882; // @[StoreQueue.scala 141:36:@827.4]
  wire  noConflicts_2; // @[StoreQueue.scala 140:95:@828.4]
  wire  _T_1885; // @[StoreQueue.scala 140:34:@830.4]
  wire  _T_1886; // @[StoreQueue.scala 140:64:@831.4]
  wire  _T_1890; // @[StoreQueue.scala 141:51:@832.4]
  wire  _T_1891; // @[StoreQueue.scala 141:36:@833.4]
  wire  noConflicts_3; // @[StoreQueue.scala 140:95:@834.4]
  wire  _T_1894; // @[StoreQueue.scala 140:34:@836.4]
  wire  _T_1895; // @[StoreQueue.scala 140:64:@837.4]
  wire  _T_1899; // @[StoreQueue.scala 141:51:@838.4]
  wire  _T_1900; // @[StoreQueue.scala 141:36:@839.4]
  wire  noConflicts_4; // @[StoreQueue.scala 140:95:@840.4]
  wire  _T_1903; // @[StoreQueue.scala 140:34:@842.4]
  wire  _T_1904; // @[StoreQueue.scala 140:64:@843.4]
  wire  _T_1908; // @[StoreQueue.scala 141:51:@844.4]
  wire  _T_1909; // @[StoreQueue.scala 141:36:@845.4]
  wire  noConflicts_5; // @[StoreQueue.scala 140:95:@846.4]
  wire  _T_1912; // @[StoreQueue.scala 140:34:@848.4]
  wire  _T_1913; // @[StoreQueue.scala 140:64:@849.4]
  wire  _T_1917; // @[StoreQueue.scala 141:51:@850.4]
  wire  _T_1918; // @[StoreQueue.scala 141:36:@851.4]
  wire  noConflicts_6; // @[StoreQueue.scala 140:95:@852.4]
  wire  _T_1921; // @[StoreQueue.scala 140:34:@854.4]
  wire  _T_1922; // @[StoreQueue.scala 140:64:@855.4]
  wire  _T_1926; // @[StoreQueue.scala 141:51:@856.4]
  wire  _T_1927; // @[StoreQueue.scala 141:36:@857.4]
  wire  noConflicts_7; // @[StoreQueue.scala 140:95:@858.4]
  wire  _GEN_265; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_266; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_267; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_268; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_269; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_270; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_271; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_273; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_274; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_275; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_276; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_277; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_278; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_279; // @[StoreQueue.scala 154:44:@860.4]
  wire  _T_1935; // @[StoreQueue.scala 154:44:@860.4]
  wire  _GEN_281; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_282; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_283; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_284; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_285; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_286; // @[StoreQueue.scala 154:66:@861.4]
  wire  _GEN_287; // @[StoreQueue.scala 154:66:@861.4]
  wire  _T_1940; // @[StoreQueue.scala 154:66:@861.4]
  wire  _T_1941; // @[StoreQueue.scala 154:63:@862.4]
  wire  _T_1944; // @[StoreQueue.scala 154:109:@864.4]
  wire  _T_1945; // @[StoreQueue.scala 154:109:@865.4]
  wire  _T_1946; // @[StoreQueue.scala 154:109:@866.4]
  wire  _T_1947; // @[StoreQueue.scala 154:109:@867.4]
  wire  _T_1948; // @[StoreQueue.scala 154:109:@868.4]
  wire  _T_1949; // @[StoreQueue.scala 154:109:@869.4]
  wire  _T_1950; // @[StoreQueue.scala 154:109:@870.4]
  wire  storeRequest; // @[StoreQueue.scala 154:88:@871.4]
  wire  _T_1953; // @[StoreQueue.scala 164:23:@876.6]
  wire  _T_1954; // @[StoreQueue.scala 164:43:@877.6]
  wire  _T_1955; // @[StoreQueue.scala 164:59:@878.6]
  wire  _GEN_288; // @[StoreQueue.scala 164:86:@879.6]
  wire  _GEN_289; // @[StoreQueue.scala 162:37:@872.4]
  wire  _T_1959; // @[StoreQueue.scala 164:23:@886.6]
  wire  _T_1960; // @[StoreQueue.scala 164:43:@887.6]
  wire  _T_1961; // @[StoreQueue.scala 164:59:@888.6]
  wire  _GEN_290; // @[StoreQueue.scala 164:86:@889.6]
  wire  _GEN_291; // @[StoreQueue.scala 162:37:@882.4]
  wire  _T_1965; // @[StoreQueue.scala 164:23:@896.6]
  wire  _T_1966; // @[StoreQueue.scala 164:43:@897.6]
  wire  _T_1967; // @[StoreQueue.scala 164:59:@898.6]
  wire  _GEN_292; // @[StoreQueue.scala 164:86:@899.6]
  wire  _GEN_293; // @[StoreQueue.scala 162:37:@892.4]
  wire  _T_1971; // @[StoreQueue.scala 164:23:@906.6]
  wire  _T_1972; // @[StoreQueue.scala 164:43:@907.6]
  wire  _T_1973; // @[StoreQueue.scala 164:59:@908.6]
  wire  _GEN_294; // @[StoreQueue.scala 164:86:@909.6]
  wire  _GEN_295; // @[StoreQueue.scala 162:37:@902.4]
  wire  _T_1977; // @[StoreQueue.scala 164:23:@916.6]
  wire  _T_1978; // @[StoreQueue.scala 164:43:@917.6]
  wire  _T_1979; // @[StoreQueue.scala 164:59:@918.6]
  wire  _GEN_296; // @[StoreQueue.scala 164:86:@919.6]
  wire  _GEN_297; // @[StoreQueue.scala 162:37:@912.4]
  wire  _T_1983; // @[StoreQueue.scala 164:23:@926.6]
  wire  _T_1984; // @[StoreQueue.scala 164:43:@927.6]
  wire  _T_1985; // @[StoreQueue.scala 164:59:@928.6]
  wire  _GEN_298; // @[StoreQueue.scala 164:86:@929.6]
  wire  _GEN_299; // @[StoreQueue.scala 162:37:@922.4]
  wire  _T_1989; // @[StoreQueue.scala 164:23:@936.6]
  wire  _T_1990; // @[StoreQueue.scala 164:43:@937.6]
  wire  _T_1991; // @[StoreQueue.scala 164:59:@938.6]
  wire  _GEN_300; // @[StoreQueue.scala 164:86:@939.6]
  wire  _GEN_301; // @[StoreQueue.scala 162:37:@932.4]
  wire  _T_1995; // @[StoreQueue.scala 164:23:@946.6]
  wire  _T_1996; // @[StoreQueue.scala 164:43:@947.6]
  wire  _T_1997; // @[StoreQueue.scala 164:59:@948.6]
  wire  _GEN_302; // @[StoreQueue.scala 164:86:@949.6]
  wire  _GEN_303; // @[StoreQueue.scala 162:37:@942.4]
  wire  entriesPorts_0_0; // @[StoreQueue.scala 180:72:@953.4]
  wire  entriesPorts_0_1; // @[StoreQueue.scala 180:72:@955.4]
  wire  entriesPorts_0_2; // @[StoreQueue.scala 180:72:@957.4]
  wire  entriesPorts_0_3; // @[StoreQueue.scala 180:72:@959.4]
  wire  entriesPorts_0_4; // @[StoreQueue.scala 180:72:@961.4]
  wire  entriesPorts_0_5; // @[StoreQueue.scala 180:72:@963.4]
  wire  entriesPorts_0_6; // @[StoreQueue.scala 180:72:@965.4]
  wire  entriesPorts_0_7; // @[StoreQueue.scala 180:72:@967.4]
  wire  _T_2410; // @[StoreQueue.scala 192:91:@987.4]
  wire  _T_2411; // @[StoreQueue.scala 192:88:@988.4]
  wire  _T_2413; // @[StoreQueue.scala 192:91:@989.4]
  wire  _T_2414; // @[StoreQueue.scala 192:88:@990.4]
  wire  _T_2416; // @[StoreQueue.scala 192:91:@991.4]
  wire  _T_2417; // @[StoreQueue.scala 192:88:@992.4]
  wire  _T_2419; // @[StoreQueue.scala 192:91:@993.4]
  wire  _T_2420; // @[StoreQueue.scala 192:88:@994.4]
  wire  _T_2422; // @[StoreQueue.scala 192:91:@995.4]
  wire  _T_2423; // @[StoreQueue.scala 192:88:@996.4]
  wire  _T_2425; // @[StoreQueue.scala 192:91:@997.4]
  wire  _T_2426; // @[StoreQueue.scala 192:88:@998.4]
  wire  _T_2428; // @[StoreQueue.scala 192:91:@999.4]
  wire  _T_2429; // @[StoreQueue.scala 192:88:@1000.4]
  wire  _T_2431; // @[StoreQueue.scala 192:91:@1001.4]
  wire  _T_2432; // @[StoreQueue.scala 192:88:@1002.4]
  wire  _T_2448; // @[StoreQueue.scala 193:91:@1012.4]
  wire  _T_2449; // @[StoreQueue.scala 193:88:@1013.4]
  wire  _T_2451; // @[StoreQueue.scala 193:91:@1014.4]
  wire  _T_2452; // @[StoreQueue.scala 193:88:@1015.4]
  wire  _T_2454; // @[StoreQueue.scala 193:91:@1016.4]
  wire  _T_2455; // @[StoreQueue.scala 193:88:@1017.4]
  wire  _T_2457; // @[StoreQueue.scala 193:91:@1018.4]
  wire  _T_2458; // @[StoreQueue.scala 193:88:@1019.4]
  wire  _T_2460; // @[StoreQueue.scala 193:91:@1020.4]
  wire  _T_2461; // @[StoreQueue.scala 193:88:@1021.4]
  wire  _T_2463; // @[StoreQueue.scala 193:91:@1022.4]
  wire  _T_2464; // @[StoreQueue.scala 193:88:@1023.4]
  wire  _T_2466; // @[StoreQueue.scala 193:91:@1024.4]
  wire  _T_2467; // @[StoreQueue.scala 193:88:@1025.4]
  wire  _T_2469; // @[StoreQueue.scala 193:91:@1026.4]
  wire  _T_2470; // @[StoreQueue.scala 193:88:@1027.4]
  wire [7:0] _T_2487; // @[OneHot.scala 52:12:@1038.4]
  wire  _T_2489; // @[util.scala 33:60:@1040.4]
  wire  _T_2490; // @[util.scala 33:60:@1041.4]
  wire  _T_2491; // @[util.scala 33:60:@1042.4]
  wire  _T_2492; // @[util.scala 33:60:@1043.4]
  wire  _T_2493; // @[util.scala 33:60:@1044.4]
  wire  _T_2494; // @[util.scala 33:60:@1045.4]
  wire  _T_2495; // @[util.scala 33:60:@1046.4]
  wire  _T_2496; // @[util.scala 33:60:@1047.4]
  wire [7:0] _T_2521; // @[Mux.scala 31:69:@1057.4]
  wire [7:0] _T_2522; // @[Mux.scala 31:69:@1058.4]
  wire [7:0] _T_2523; // @[Mux.scala 31:69:@1059.4]
  wire [7:0] _T_2524; // @[Mux.scala 31:69:@1060.4]
  wire [7:0] _T_2525; // @[Mux.scala 31:69:@1061.4]
  wire [7:0] _T_2526; // @[Mux.scala 31:69:@1062.4]
  wire [7:0] _T_2527; // @[Mux.scala 31:69:@1063.4]
  wire [7:0] _T_2528; // @[Mux.scala 31:69:@1064.4]
  wire  _T_2529; // @[OneHot.scala 66:30:@1065.4]
  wire  _T_2530; // @[OneHot.scala 66:30:@1066.4]
  wire  _T_2531; // @[OneHot.scala 66:30:@1067.4]
  wire  _T_2532; // @[OneHot.scala 66:30:@1068.4]
  wire  _T_2533; // @[OneHot.scala 66:30:@1069.4]
  wire  _T_2534; // @[OneHot.scala 66:30:@1070.4]
  wire  _T_2535; // @[OneHot.scala 66:30:@1071.4]
  wire  _T_2536; // @[OneHot.scala 66:30:@1072.4]
  wire [7:0] _T_2561; // @[Mux.scala 31:69:@1082.4]
  wire [7:0] _T_2562; // @[Mux.scala 31:69:@1083.4]
  wire [7:0] _T_2563; // @[Mux.scala 31:69:@1084.4]
  wire [7:0] _T_2564; // @[Mux.scala 31:69:@1085.4]
  wire [7:0] _T_2565; // @[Mux.scala 31:69:@1086.4]
  wire [7:0] _T_2566; // @[Mux.scala 31:69:@1087.4]
  wire [7:0] _T_2567; // @[Mux.scala 31:69:@1088.4]
  wire [7:0] _T_2568; // @[Mux.scala 31:69:@1089.4]
  wire  _T_2569; // @[OneHot.scala 66:30:@1090.4]
  wire  _T_2570; // @[OneHot.scala 66:30:@1091.4]
  wire  _T_2571; // @[OneHot.scala 66:30:@1092.4]
  wire  _T_2572; // @[OneHot.scala 66:30:@1093.4]
  wire  _T_2573; // @[OneHot.scala 66:30:@1094.4]
  wire  _T_2574; // @[OneHot.scala 66:30:@1095.4]
  wire  _T_2575; // @[OneHot.scala 66:30:@1096.4]
  wire  _T_2576; // @[OneHot.scala 66:30:@1097.4]
  wire [7:0] _T_2601; // @[Mux.scala 31:69:@1107.4]
  wire [7:0] _T_2602; // @[Mux.scala 31:69:@1108.4]
  wire [7:0] _T_2603; // @[Mux.scala 31:69:@1109.4]
  wire [7:0] _T_2604; // @[Mux.scala 31:69:@1110.4]
  wire [7:0] _T_2605; // @[Mux.scala 31:69:@1111.4]
  wire [7:0] _T_2606; // @[Mux.scala 31:69:@1112.4]
  wire [7:0] _T_2607; // @[Mux.scala 31:69:@1113.4]
  wire [7:0] _T_2608; // @[Mux.scala 31:69:@1114.4]
  wire  _T_2609; // @[OneHot.scala 66:30:@1115.4]
  wire  _T_2610; // @[OneHot.scala 66:30:@1116.4]
  wire  _T_2611; // @[OneHot.scala 66:30:@1117.4]
  wire  _T_2612; // @[OneHot.scala 66:30:@1118.4]
  wire  _T_2613; // @[OneHot.scala 66:30:@1119.4]
  wire  _T_2614; // @[OneHot.scala 66:30:@1120.4]
  wire  _T_2615; // @[OneHot.scala 66:30:@1121.4]
  wire  _T_2616; // @[OneHot.scala 66:30:@1122.4]
  wire [7:0] _T_2641; // @[Mux.scala 31:69:@1132.4]
  wire [7:0] _T_2642; // @[Mux.scala 31:69:@1133.4]
  wire [7:0] _T_2643; // @[Mux.scala 31:69:@1134.4]
  wire [7:0] _T_2644; // @[Mux.scala 31:69:@1135.4]
  wire [7:0] _T_2645; // @[Mux.scala 31:69:@1136.4]
  wire [7:0] _T_2646; // @[Mux.scala 31:69:@1137.4]
  wire [7:0] _T_2647; // @[Mux.scala 31:69:@1138.4]
  wire [7:0] _T_2648; // @[Mux.scala 31:69:@1139.4]
  wire  _T_2649; // @[OneHot.scala 66:30:@1140.4]
  wire  _T_2650; // @[OneHot.scala 66:30:@1141.4]
  wire  _T_2651; // @[OneHot.scala 66:30:@1142.4]
  wire  _T_2652; // @[OneHot.scala 66:30:@1143.4]
  wire  _T_2653; // @[OneHot.scala 66:30:@1144.4]
  wire  _T_2654; // @[OneHot.scala 66:30:@1145.4]
  wire  _T_2655; // @[OneHot.scala 66:30:@1146.4]
  wire  _T_2656; // @[OneHot.scala 66:30:@1147.4]
  wire [7:0] _T_2681; // @[Mux.scala 31:69:@1157.4]
  wire [7:0] _T_2682; // @[Mux.scala 31:69:@1158.4]
  wire [7:0] _T_2683; // @[Mux.scala 31:69:@1159.4]
  wire [7:0] _T_2684; // @[Mux.scala 31:69:@1160.4]
  wire [7:0] _T_2685; // @[Mux.scala 31:69:@1161.4]
  wire [7:0] _T_2686; // @[Mux.scala 31:69:@1162.4]
  wire [7:0] _T_2687; // @[Mux.scala 31:69:@1163.4]
  wire [7:0] _T_2688; // @[Mux.scala 31:69:@1164.4]
  wire  _T_2689; // @[OneHot.scala 66:30:@1165.4]
  wire  _T_2690; // @[OneHot.scala 66:30:@1166.4]
  wire  _T_2691; // @[OneHot.scala 66:30:@1167.4]
  wire  _T_2692; // @[OneHot.scala 66:30:@1168.4]
  wire  _T_2693; // @[OneHot.scala 66:30:@1169.4]
  wire  _T_2694; // @[OneHot.scala 66:30:@1170.4]
  wire  _T_2695; // @[OneHot.scala 66:30:@1171.4]
  wire  _T_2696; // @[OneHot.scala 66:30:@1172.4]
  wire [7:0] _T_2721; // @[Mux.scala 31:69:@1182.4]
  wire [7:0] _T_2722; // @[Mux.scala 31:69:@1183.4]
  wire [7:0] _T_2723; // @[Mux.scala 31:69:@1184.4]
  wire [7:0] _T_2724; // @[Mux.scala 31:69:@1185.4]
  wire [7:0] _T_2725; // @[Mux.scala 31:69:@1186.4]
  wire [7:0] _T_2726; // @[Mux.scala 31:69:@1187.4]
  wire [7:0] _T_2727; // @[Mux.scala 31:69:@1188.4]
  wire [7:0] _T_2728; // @[Mux.scala 31:69:@1189.4]
  wire  _T_2729; // @[OneHot.scala 66:30:@1190.4]
  wire  _T_2730; // @[OneHot.scala 66:30:@1191.4]
  wire  _T_2731; // @[OneHot.scala 66:30:@1192.4]
  wire  _T_2732; // @[OneHot.scala 66:30:@1193.4]
  wire  _T_2733; // @[OneHot.scala 66:30:@1194.4]
  wire  _T_2734; // @[OneHot.scala 66:30:@1195.4]
  wire  _T_2735; // @[OneHot.scala 66:30:@1196.4]
  wire  _T_2736; // @[OneHot.scala 66:30:@1197.4]
  wire [7:0] _T_2761; // @[Mux.scala 31:69:@1207.4]
  wire [7:0] _T_2762; // @[Mux.scala 31:69:@1208.4]
  wire [7:0] _T_2763; // @[Mux.scala 31:69:@1209.4]
  wire [7:0] _T_2764; // @[Mux.scala 31:69:@1210.4]
  wire [7:0] _T_2765; // @[Mux.scala 31:69:@1211.4]
  wire [7:0] _T_2766; // @[Mux.scala 31:69:@1212.4]
  wire [7:0] _T_2767; // @[Mux.scala 31:69:@1213.4]
  wire [7:0] _T_2768; // @[Mux.scala 31:69:@1214.4]
  wire  _T_2769; // @[OneHot.scala 66:30:@1215.4]
  wire  _T_2770; // @[OneHot.scala 66:30:@1216.4]
  wire  _T_2771; // @[OneHot.scala 66:30:@1217.4]
  wire  _T_2772; // @[OneHot.scala 66:30:@1218.4]
  wire  _T_2773; // @[OneHot.scala 66:30:@1219.4]
  wire  _T_2774; // @[OneHot.scala 66:30:@1220.4]
  wire  _T_2775; // @[OneHot.scala 66:30:@1221.4]
  wire  _T_2776; // @[OneHot.scala 66:30:@1222.4]
  wire [7:0] _T_2801; // @[Mux.scala 31:69:@1232.4]
  wire [7:0] _T_2802; // @[Mux.scala 31:69:@1233.4]
  wire [7:0] _T_2803; // @[Mux.scala 31:69:@1234.4]
  wire [7:0] _T_2804; // @[Mux.scala 31:69:@1235.4]
  wire [7:0] _T_2805; // @[Mux.scala 31:69:@1236.4]
  wire [7:0] _T_2806; // @[Mux.scala 31:69:@1237.4]
  wire [7:0] _T_2807; // @[Mux.scala 31:69:@1238.4]
  wire [7:0] _T_2808; // @[Mux.scala 31:69:@1239.4]
  wire  _T_2809; // @[OneHot.scala 66:30:@1240.4]
  wire  _T_2810; // @[OneHot.scala 66:30:@1241.4]
  wire  _T_2811; // @[OneHot.scala 66:30:@1242.4]
  wire  _T_2812; // @[OneHot.scala 66:30:@1243.4]
  wire  _T_2813; // @[OneHot.scala 66:30:@1244.4]
  wire  _T_2814; // @[OneHot.scala 66:30:@1245.4]
  wire  _T_2815; // @[OneHot.scala 66:30:@1246.4]
  wire  _T_2816; // @[OneHot.scala 66:30:@1247.4]
  wire [7:0] _T_2857; // @[Mux.scala 19:72:@1263.4]
  wire [7:0] _T_2859; // @[Mux.scala 19:72:@1264.4]
  wire [7:0] _T_2866; // @[Mux.scala 19:72:@1271.4]
  wire [7:0] _T_2868; // @[Mux.scala 19:72:@1272.4]
  wire [7:0] _T_2875; // @[Mux.scala 19:72:@1279.4]
  wire [7:0] _T_2877; // @[Mux.scala 19:72:@1280.4]
  wire [7:0] _T_2884; // @[Mux.scala 19:72:@1287.4]
  wire [7:0] _T_2886; // @[Mux.scala 19:72:@1288.4]
  wire [7:0] _T_2893; // @[Mux.scala 19:72:@1295.4]
  wire [7:0] _T_2895; // @[Mux.scala 19:72:@1296.4]
  wire [7:0] _T_2902; // @[Mux.scala 19:72:@1303.4]
  wire [7:0] _T_2904; // @[Mux.scala 19:72:@1304.4]
  wire [7:0] _T_2911; // @[Mux.scala 19:72:@1311.4]
  wire [7:0] _T_2913; // @[Mux.scala 19:72:@1312.4]
  wire [7:0] _T_2920; // @[Mux.scala 19:72:@1319.4]
  wire [7:0] _T_2922; // @[Mux.scala 19:72:@1320.4]
  wire [7:0] _T_2923; // @[Mux.scala 19:72:@1321.4]
  wire [7:0] _T_2924; // @[Mux.scala 19:72:@1322.4]
  wire [7:0] _T_2925; // @[Mux.scala 19:72:@1323.4]
  wire [7:0] _T_2926; // @[Mux.scala 19:72:@1324.4]
  wire [7:0] _T_2927; // @[Mux.scala 19:72:@1325.4]
  wire [7:0] _T_2928; // @[Mux.scala 19:72:@1326.4]
  wire [7:0] _T_2929; // @[Mux.scala 19:72:@1327.4]
  wire  inputAddrPriorityPorts_0_0; // @[Mux.scala 19:72:@1331.4]
  wire  inputAddrPriorityPorts_0_1; // @[Mux.scala 19:72:@1333.4]
  wire  inputAddrPriorityPorts_0_2; // @[Mux.scala 19:72:@1335.4]
  wire  inputAddrPriorityPorts_0_3; // @[Mux.scala 19:72:@1337.4]
  wire  inputAddrPriorityPorts_0_4; // @[Mux.scala 19:72:@1339.4]
  wire  inputAddrPriorityPorts_0_5; // @[Mux.scala 19:72:@1341.4]
  wire  inputAddrPriorityPorts_0_6; // @[Mux.scala 19:72:@1343.4]
  wire  inputAddrPriorityPorts_0_7; // @[Mux.scala 19:72:@1345.4]
  wire [7:0] _T_3043; // @[Mux.scala 31:69:@1375.4]
  wire [7:0] _T_3044; // @[Mux.scala 31:69:@1376.4]
  wire [7:0] _T_3045; // @[Mux.scala 31:69:@1377.4]
  wire [7:0] _T_3046; // @[Mux.scala 31:69:@1378.4]
  wire [7:0] _T_3047; // @[Mux.scala 31:69:@1379.4]
  wire [7:0] _T_3048; // @[Mux.scala 31:69:@1380.4]
  wire [7:0] _T_3049; // @[Mux.scala 31:69:@1381.4]
  wire [7:0] _T_3050; // @[Mux.scala 31:69:@1382.4]
  wire  _T_3051; // @[OneHot.scala 66:30:@1383.4]
  wire  _T_3052; // @[OneHot.scala 66:30:@1384.4]
  wire  _T_3053; // @[OneHot.scala 66:30:@1385.4]
  wire  _T_3054; // @[OneHot.scala 66:30:@1386.4]
  wire  _T_3055; // @[OneHot.scala 66:30:@1387.4]
  wire  _T_3056; // @[OneHot.scala 66:30:@1388.4]
  wire  _T_3057; // @[OneHot.scala 66:30:@1389.4]
  wire  _T_3058; // @[OneHot.scala 66:30:@1390.4]
  wire [7:0] _T_3083; // @[Mux.scala 31:69:@1400.4]
  wire [7:0] _T_3084; // @[Mux.scala 31:69:@1401.4]
  wire [7:0] _T_3085; // @[Mux.scala 31:69:@1402.4]
  wire [7:0] _T_3086; // @[Mux.scala 31:69:@1403.4]
  wire [7:0] _T_3087; // @[Mux.scala 31:69:@1404.4]
  wire [7:0] _T_3088; // @[Mux.scala 31:69:@1405.4]
  wire [7:0] _T_3089; // @[Mux.scala 31:69:@1406.4]
  wire [7:0] _T_3090; // @[Mux.scala 31:69:@1407.4]
  wire  _T_3091; // @[OneHot.scala 66:30:@1408.4]
  wire  _T_3092; // @[OneHot.scala 66:30:@1409.4]
  wire  _T_3093; // @[OneHot.scala 66:30:@1410.4]
  wire  _T_3094; // @[OneHot.scala 66:30:@1411.4]
  wire  _T_3095; // @[OneHot.scala 66:30:@1412.4]
  wire  _T_3096; // @[OneHot.scala 66:30:@1413.4]
  wire  _T_3097; // @[OneHot.scala 66:30:@1414.4]
  wire  _T_3098; // @[OneHot.scala 66:30:@1415.4]
  wire [7:0] _T_3123; // @[Mux.scala 31:69:@1425.4]
  wire [7:0] _T_3124; // @[Mux.scala 31:69:@1426.4]
  wire [7:0] _T_3125; // @[Mux.scala 31:69:@1427.4]
  wire [7:0] _T_3126; // @[Mux.scala 31:69:@1428.4]
  wire [7:0] _T_3127; // @[Mux.scala 31:69:@1429.4]
  wire [7:0] _T_3128; // @[Mux.scala 31:69:@1430.4]
  wire [7:0] _T_3129; // @[Mux.scala 31:69:@1431.4]
  wire [7:0] _T_3130; // @[Mux.scala 31:69:@1432.4]
  wire  _T_3131; // @[OneHot.scala 66:30:@1433.4]
  wire  _T_3132; // @[OneHot.scala 66:30:@1434.4]
  wire  _T_3133; // @[OneHot.scala 66:30:@1435.4]
  wire  _T_3134; // @[OneHot.scala 66:30:@1436.4]
  wire  _T_3135; // @[OneHot.scala 66:30:@1437.4]
  wire  _T_3136; // @[OneHot.scala 66:30:@1438.4]
  wire  _T_3137; // @[OneHot.scala 66:30:@1439.4]
  wire  _T_3138; // @[OneHot.scala 66:30:@1440.4]
  wire [7:0] _T_3163; // @[Mux.scala 31:69:@1450.4]
  wire [7:0] _T_3164; // @[Mux.scala 31:69:@1451.4]
  wire [7:0] _T_3165; // @[Mux.scala 31:69:@1452.4]
  wire [7:0] _T_3166; // @[Mux.scala 31:69:@1453.4]
  wire [7:0] _T_3167; // @[Mux.scala 31:69:@1454.4]
  wire [7:0] _T_3168; // @[Mux.scala 31:69:@1455.4]
  wire [7:0] _T_3169; // @[Mux.scala 31:69:@1456.4]
  wire [7:0] _T_3170; // @[Mux.scala 31:69:@1457.4]
  wire  _T_3171; // @[OneHot.scala 66:30:@1458.4]
  wire  _T_3172; // @[OneHot.scala 66:30:@1459.4]
  wire  _T_3173; // @[OneHot.scala 66:30:@1460.4]
  wire  _T_3174; // @[OneHot.scala 66:30:@1461.4]
  wire  _T_3175; // @[OneHot.scala 66:30:@1462.4]
  wire  _T_3176; // @[OneHot.scala 66:30:@1463.4]
  wire  _T_3177; // @[OneHot.scala 66:30:@1464.4]
  wire  _T_3178; // @[OneHot.scala 66:30:@1465.4]
  wire [7:0] _T_3203; // @[Mux.scala 31:69:@1475.4]
  wire [7:0] _T_3204; // @[Mux.scala 31:69:@1476.4]
  wire [7:0] _T_3205; // @[Mux.scala 31:69:@1477.4]
  wire [7:0] _T_3206; // @[Mux.scala 31:69:@1478.4]
  wire [7:0] _T_3207; // @[Mux.scala 31:69:@1479.4]
  wire [7:0] _T_3208; // @[Mux.scala 31:69:@1480.4]
  wire [7:0] _T_3209; // @[Mux.scala 31:69:@1481.4]
  wire [7:0] _T_3210; // @[Mux.scala 31:69:@1482.4]
  wire  _T_3211; // @[OneHot.scala 66:30:@1483.4]
  wire  _T_3212; // @[OneHot.scala 66:30:@1484.4]
  wire  _T_3213; // @[OneHot.scala 66:30:@1485.4]
  wire  _T_3214; // @[OneHot.scala 66:30:@1486.4]
  wire  _T_3215; // @[OneHot.scala 66:30:@1487.4]
  wire  _T_3216; // @[OneHot.scala 66:30:@1488.4]
  wire  _T_3217; // @[OneHot.scala 66:30:@1489.4]
  wire  _T_3218; // @[OneHot.scala 66:30:@1490.4]
  wire [7:0] _T_3243; // @[Mux.scala 31:69:@1500.4]
  wire [7:0] _T_3244; // @[Mux.scala 31:69:@1501.4]
  wire [7:0] _T_3245; // @[Mux.scala 31:69:@1502.4]
  wire [7:0] _T_3246; // @[Mux.scala 31:69:@1503.4]
  wire [7:0] _T_3247; // @[Mux.scala 31:69:@1504.4]
  wire [7:0] _T_3248; // @[Mux.scala 31:69:@1505.4]
  wire [7:0] _T_3249; // @[Mux.scala 31:69:@1506.4]
  wire [7:0] _T_3250; // @[Mux.scala 31:69:@1507.4]
  wire  _T_3251; // @[OneHot.scala 66:30:@1508.4]
  wire  _T_3252; // @[OneHot.scala 66:30:@1509.4]
  wire  _T_3253; // @[OneHot.scala 66:30:@1510.4]
  wire  _T_3254; // @[OneHot.scala 66:30:@1511.4]
  wire  _T_3255; // @[OneHot.scala 66:30:@1512.4]
  wire  _T_3256; // @[OneHot.scala 66:30:@1513.4]
  wire  _T_3257; // @[OneHot.scala 66:30:@1514.4]
  wire  _T_3258; // @[OneHot.scala 66:30:@1515.4]
  wire [7:0] _T_3283; // @[Mux.scala 31:69:@1525.4]
  wire [7:0] _T_3284; // @[Mux.scala 31:69:@1526.4]
  wire [7:0] _T_3285; // @[Mux.scala 31:69:@1527.4]
  wire [7:0] _T_3286; // @[Mux.scala 31:69:@1528.4]
  wire [7:0] _T_3287; // @[Mux.scala 31:69:@1529.4]
  wire [7:0] _T_3288; // @[Mux.scala 31:69:@1530.4]
  wire [7:0] _T_3289; // @[Mux.scala 31:69:@1531.4]
  wire [7:0] _T_3290; // @[Mux.scala 31:69:@1532.4]
  wire  _T_3291; // @[OneHot.scala 66:30:@1533.4]
  wire  _T_3292; // @[OneHot.scala 66:30:@1534.4]
  wire  _T_3293; // @[OneHot.scala 66:30:@1535.4]
  wire  _T_3294; // @[OneHot.scala 66:30:@1536.4]
  wire  _T_3295; // @[OneHot.scala 66:30:@1537.4]
  wire  _T_3296; // @[OneHot.scala 66:30:@1538.4]
  wire  _T_3297; // @[OneHot.scala 66:30:@1539.4]
  wire  _T_3298; // @[OneHot.scala 66:30:@1540.4]
  wire [7:0] _T_3323; // @[Mux.scala 31:69:@1550.4]
  wire [7:0] _T_3324; // @[Mux.scala 31:69:@1551.4]
  wire [7:0] _T_3325; // @[Mux.scala 31:69:@1552.4]
  wire [7:0] _T_3326; // @[Mux.scala 31:69:@1553.4]
  wire [7:0] _T_3327; // @[Mux.scala 31:69:@1554.4]
  wire [7:0] _T_3328; // @[Mux.scala 31:69:@1555.4]
  wire [7:0] _T_3329; // @[Mux.scala 31:69:@1556.4]
  wire [7:0] _T_3330; // @[Mux.scala 31:69:@1557.4]
  wire  _T_3331; // @[OneHot.scala 66:30:@1558.4]
  wire  _T_3332; // @[OneHot.scala 66:30:@1559.4]
  wire  _T_3333; // @[OneHot.scala 66:30:@1560.4]
  wire  _T_3334; // @[OneHot.scala 66:30:@1561.4]
  wire  _T_3335; // @[OneHot.scala 66:30:@1562.4]
  wire  _T_3336; // @[OneHot.scala 66:30:@1563.4]
  wire  _T_3337; // @[OneHot.scala 66:30:@1564.4]
  wire  _T_3338; // @[OneHot.scala 66:30:@1565.4]
  wire [7:0] _T_3379; // @[Mux.scala 19:72:@1581.4]
  wire [7:0] _T_3381; // @[Mux.scala 19:72:@1582.4]
  wire [7:0] _T_3388; // @[Mux.scala 19:72:@1589.4]
  wire [7:0] _T_3390; // @[Mux.scala 19:72:@1590.4]
  wire [7:0] _T_3397; // @[Mux.scala 19:72:@1597.4]
  wire [7:0] _T_3399; // @[Mux.scala 19:72:@1598.4]
  wire [7:0] _T_3406; // @[Mux.scala 19:72:@1605.4]
  wire [7:0] _T_3408; // @[Mux.scala 19:72:@1606.4]
  wire [7:0] _T_3415; // @[Mux.scala 19:72:@1613.4]
  wire [7:0] _T_3417; // @[Mux.scala 19:72:@1614.4]
  wire [7:0] _T_3424; // @[Mux.scala 19:72:@1621.4]
  wire [7:0] _T_3426; // @[Mux.scala 19:72:@1622.4]
  wire [7:0] _T_3433; // @[Mux.scala 19:72:@1629.4]
  wire [7:0] _T_3435; // @[Mux.scala 19:72:@1630.4]
  wire [7:0] _T_3442; // @[Mux.scala 19:72:@1637.4]
  wire [7:0] _T_3444; // @[Mux.scala 19:72:@1638.4]
  wire [7:0] _T_3445; // @[Mux.scala 19:72:@1639.4]
  wire [7:0] _T_3446; // @[Mux.scala 19:72:@1640.4]
  wire [7:0] _T_3447; // @[Mux.scala 19:72:@1641.4]
  wire [7:0] _T_3448; // @[Mux.scala 19:72:@1642.4]
  wire [7:0] _T_3449; // @[Mux.scala 19:72:@1643.4]
  wire [7:0] _T_3450; // @[Mux.scala 19:72:@1644.4]
  wire [7:0] _T_3451; // @[Mux.scala 19:72:@1645.4]
  wire  inputDataPriorityPorts_0_0; // @[Mux.scala 19:72:@1649.4]
  wire  inputDataPriorityPorts_0_1; // @[Mux.scala 19:72:@1651.4]
  wire  inputDataPriorityPorts_0_2; // @[Mux.scala 19:72:@1653.4]
  wire  inputDataPriorityPorts_0_3; // @[Mux.scala 19:72:@1655.4]
  wire  inputDataPriorityPorts_0_4; // @[Mux.scala 19:72:@1657.4]
  wire  inputDataPriorityPorts_0_5; // @[Mux.scala 19:72:@1659.4]
  wire  inputDataPriorityPorts_0_6; // @[Mux.scala 19:72:@1661.4]
  wire  inputDataPriorityPorts_0_7; // @[Mux.scala 19:72:@1663.4]
  wire  _T_3531; // @[StoreQueue.scala 192:88:@1674.4]
  wire  _T_3534; // @[StoreQueue.scala 192:88:@1676.4]
  wire  _T_3537; // @[StoreQueue.scala 192:88:@1678.4]
  wire  _T_3540; // @[StoreQueue.scala 192:88:@1680.4]
  wire  _T_3543; // @[StoreQueue.scala 192:88:@1682.4]
  wire  _T_3546; // @[StoreQueue.scala 192:88:@1684.4]
  wire  _T_3549; // @[StoreQueue.scala 192:88:@1686.4]
  wire  _T_3552; // @[StoreQueue.scala 192:88:@1688.4]
  wire  _T_3569; // @[StoreQueue.scala 193:88:@1699.4]
  wire  _T_3572; // @[StoreQueue.scala 193:88:@1701.4]
  wire  _T_3575; // @[StoreQueue.scala 193:88:@1703.4]
  wire  _T_3578; // @[StoreQueue.scala 193:88:@1705.4]
  wire  _T_3581; // @[StoreQueue.scala 193:88:@1707.4]
  wire  _T_3584; // @[StoreQueue.scala 193:88:@1709.4]
  wire  _T_3587; // @[StoreQueue.scala 193:88:@1711.4]
  wire  _T_3590; // @[StoreQueue.scala 193:88:@1713.4]
  wire [7:0] _T_3641; // @[Mux.scala 31:69:@1743.4]
  wire [7:0] _T_3642; // @[Mux.scala 31:69:@1744.4]
  wire [7:0] _T_3643; // @[Mux.scala 31:69:@1745.4]
  wire [7:0] _T_3644; // @[Mux.scala 31:69:@1746.4]
  wire [7:0] _T_3645; // @[Mux.scala 31:69:@1747.4]
  wire [7:0] _T_3646; // @[Mux.scala 31:69:@1748.4]
  wire [7:0] _T_3647; // @[Mux.scala 31:69:@1749.4]
  wire [7:0] _T_3648; // @[Mux.scala 31:69:@1750.4]
  wire  _T_3649; // @[OneHot.scala 66:30:@1751.4]
  wire  _T_3650; // @[OneHot.scala 66:30:@1752.4]
  wire  _T_3651; // @[OneHot.scala 66:30:@1753.4]
  wire  _T_3652; // @[OneHot.scala 66:30:@1754.4]
  wire  _T_3653; // @[OneHot.scala 66:30:@1755.4]
  wire  _T_3654; // @[OneHot.scala 66:30:@1756.4]
  wire  _T_3655; // @[OneHot.scala 66:30:@1757.4]
  wire  _T_3656; // @[OneHot.scala 66:30:@1758.4]
  wire [7:0] _T_3681; // @[Mux.scala 31:69:@1768.4]
  wire [7:0] _T_3682; // @[Mux.scala 31:69:@1769.4]
  wire [7:0] _T_3683; // @[Mux.scala 31:69:@1770.4]
  wire [7:0] _T_3684; // @[Mux.scala 31:69:@1771.4]
  wire [7:0] _T_3685; // @[Mux.scala 31:69:@1772.4]
  wire [7:0] _T_3686; // @[Mux.scala 31:69:@1773.4]
  wire [7:0] _T_3687; // @[Mux.scala 31:69:@1774.4]
  wire [7:0] _T_3688; // @[Mux.scala 31:69:@1775.4]
  wire  _T_3689; // @[OneHot.scala 66:30:@1776.4]
  wire  _T_3690; // @[OneHot.scala 66:30:@1777.4]
  wire  _T_3691; // @[OneHot.scala 66:30:@1778.4]
  wire  _T_3692; // @[OneHot.scala 66:30:@1779.4]
  wire  _T_3693; // @[OneHot.scala 66:30:@1780.4]
  wire  _T_3694; // @[OneHot.scala 66:30:@1781.4]
  wire  _T_3695; // @[OneHot.scala 66:30:@1782.4]
  wire  _T_3696; // @[OneHot.scala 66:30:@1783.4]
  wire [7:0] _T_3721; // @[Mux.scala 31:69:@1793.4]
  wire [7:0] _T_3722; // @[Mux.scala 31:69:@1794.4]
  wire [7:0] _T_3723; // @[Mux.scala 31:69:@1795.4]
  wire [7:0] _T_3724; // @[Mux.scala 31:69:@1796.4]
  wire [7:0] _T_3725; // @[Mux.scala 31:69:@1797.4]
  wire [7:0] _T_3726; // @[Mux.scala 31:69:@1798.4]
  wire [7:0] _T_3727; // @[Mux.scala 31:69:@1799.4]
  wire [7:0] _T_3728; // @[Mux.scala 31:69:@1800.4]
  wire  _T_3729; // @[OneHot.scala 66:30:@1801.4]
  wire  _T_3730; // @[OneHot.scala 66:30:@1802.4]
  wire  _T_3731; // @[OneHot.scala 66:30:@1803.4]
  wire  _T_3732; // @[OneHot.scala 66:30:@1804.4]
  wire  _T_3733; // @[OneHot.scala 66:30:@1805.4]
  wire  _T_3734; // @[OneHot.scala 66:30:@1806.4]
  wire  _T_3735; // @[OneHot.scala 66:30:@1807.4]
  wire  _T_3736; // @[OneHot.scala 66:30:@1808.4]
  wire [7:0] _T_3761; // @[Mux.scala 31:69:@1818.4]
  wire [7:0] _T_3762; // @[Mux.scala 31:69:@1819.4]
  wire [7:0] _T_3763; // @[Mux.scala 31:69:@1820.4]
  wire [7:0] _T_3764; // @[Mux.scala 31:69:@1821.4]
  wire [7:0] _T_3765; // @[Mux.scala 31:69:@1822.4]
  wire [7:0] _T_3766; // @[Mux.scala 31:69:@1823.4]
  wire [7:0] _T_3767; // @[Mux.scala 31:69:@1824.4]
  wire [7:0] _T_3768; // @[Mux.scala 31:69:@1825.4]
  wire  _T_3769; // @[OneHot.scala 66:30:@1826.4]
  wire  _T_3770; // @[OneHot.scala 66:30:@1827.4]
  wire  _T_3771; // @[OneHot.scala 66:30:@1828.4]
  wire  _T_3772; // @[OneHot.scala 66:30:@1829.4]
  wire  _T_3773; // @[OneHot.scala 66:30:@1830.4]
  wire  _T_3774; // @[OneHot.scala 66:30:@1831.4]
  wire  _T_3775; // @[OneHot.scala 66:30:@1832.4]
  wire  _T_3776; // @[OneHot.scala 66:30:@1833.4]
  wire [7:0] _T_3801; // @[Mux.scala 31:69:@1843.4]
  wire [7:0] _T_3802; // @[Mux.scala 31:69:@1844.4]
  wire [7:0] _T_3803; // @[Mux.scala 31:69:@1845.4]
  wire [7:0] _T_3804; // @[Mux.scala 31:69:@1846.4]
  wire [7:0] _T_3805; // @[Mux.scala 31:69:@1847.4]
  wire [7:0] _T_3806; // @[Mux.scala 31:69:@1848.4]
  wire [7:0] _T_3807; // @[Mux.scala 31:69:@1849.4]
  wire [7:0] _T_3808; // @[Mux.scala 31:69:@1850.4]
  wire  _T_3809; // @[OneHot.scala 66:30:@1851.4]
  wire  _T_3810; // @[OneHot.scala 66:30:@1852.4]
  wire  _T_3811; // @[OneHot.scala 66:30:@1853.4]
  wire  _T_3812; // @[OneHot.scala 66:30:@1854.4]
  wire  _T_3813; // @[OneHot.scala 66:30:@1855.4]
  wire  _T_3814; // @[OneHot.scala 66:30:@1856.4]
  wire  _T_3815; // @[OneHot.scala 66:30:@1857.4]
  wire  _T_3816; // @[OneHot.scala 66:30:@1858.4]
  wire [7:0] _T_3841; // @[Mux.scala 31:69:@1868.4]
  wire [7:0] _T_3842; // @[Mux.scala 31:69:@1869.4]
  wire [7:0] _T_3843; // @[Mux.scala 31:69:@1870.4]
  wire [7:0] _T_3844; // @[Mux.scala 31:69:@1871.4]
  wire [7:0] _T_3845; // @[Mux.scala 31:69:@1872.4]
  wire [7:0] _T_3846; // @[Mux.scala 31:69:@1873.4]
  wire [7:0] _T_3847; // @[Mux.scala 31:69:@1874.4]
  wire [7:0] _T_3848; // @[Mux.scala 31:69:@1875.4]
  wire  _T_3849; // @[OneHot.scala 66:30:@1876.4]
  wire  _T_3850; // @[OneHot.scala 66:30:@1877.4]
  wire  _T_3851; // @[OneHot.scala 66:30:@1878.4]
  wire  _T_3852; // @[OneHot.scala 66:30:@1879.4]
  wire  _T_3853; // @[OneHot.scala 66:30:@1880.4]
  wire  _T_3854; // @[OneHot.scala 66:30:@1881.4]
  wire  _T_3855; // @[OneHot.scala 66:30:@1882.4]
  wire  _T_3856; // @[OneHot.scala 66:30:@1883.4]
  wire [7:0] _T_3881; // @[Mux.scala 31:69:@1893.4]
  wire [7:0] _T_3882; // @[Mux.scala 31:69:@1894.4]
  wire [7:0] _T_3883; // @[Mux.scala 31:69:@1895.4]
  wire [7:0] _T_3884; // @[Mux.scala 31:69:@1896.4]
  wire [7:0] _T_3885; // @[Mux.scala 31:69:@1897.4]
  wire [7:0] _T_3886; // @[Mux.scala 31:69:@1898.4]
  wire [7:0] _T_3887; // @[Mux.scala 31:69:@1899.4]
  wire [7:0] _T_3888; // @[Mux.scala 31:69:@1900.4]
  wire  _T_3889; // @[OneHot.scala 66:30:@1901.4]
  wire  _T_3890; // @[OneHot.scala 66:30:@1902.4]
  wire  _T_3891; // @[OneHot.scala 66:30:@1903.4]
  wire  _T_3892; // @[OneHot.scala 66:30:@1904.4]
  wire  _T_3893; // @[OneHot.scala 66:30:@1905.4]
  wire  _T_3894; // @[OneHot.scala 66:30:@1906.4]
  wire  _T_3895; // @[OneHot.scala 66:30:@1907.4]
  wire  _T_3896; // @[OneHot.scala 66:30:@1908.4]
  wire [7:0] _T_3921; // @[Mux.scala 31:69:@1918.4]
  wire [7:0] _T_3922; // @[Mux.scala 31:69:@1919.4]
  wire [7:0] _T_3923; // @[Mux.scala 31:69:@1920.4]
  wire [7:0] _T_3924; // @[Mux.scala 31:69:@1921.4]
  wire [7:0] _T_3925; // @[Mux.scala 31:69:@1922.4]
  wire [7:0] _T_3926; // @[Mux.scala 31:69:@1923.4]
  wire [7:0] _T_3927; // @[Mux.scala 31:69:@1924.4]
  wire [7:0] _T_3928; // @[Mux.scala 31:69:@1925.4]
  wire  _T_3929; // @[OneHot.scala 66:30:@1926.4]
  wire  _T_3930; // @[OneHot.scala 66:30:@1927.4]
  wire  _T_3931; // @[OneHot.scala 66:30:@1928.4]
  wire  _T_3932; // @[OneHot.scala 66:30:@1929.4]
  wire  _T_3933; // @[OneHot.scala 66:30:@1930.4]
  wire  _T_3934; // @[OneHot.scala 66:30:@1931.4]
  wire  _T_3935; // @[OneHot.scala 66:30:@1932.4]
  wire  _T_3936; // @[OneHot.scala 66:30:@1933.4]
  wire [7:0] _T_3977; // @[Mux.scala 19:72:@1949.4]
  wire [7:0] _T_3979; // @[Mux.scala 19:72:@1950.4]
  wire [7:0] _T_3986; // @[Mux.scala 19:72:@1957.4]
  wire [7:0] _T_3988; // @[Mux.scala 19:72:@1958.4]
  wire [7:0] _T_3995; // @[Mux.scala 19:72:@1965.4]
  wire [7:0] _T_3997; // @[Mux.scala 19:72:@1966.4]
  wire [7:0] _T_4004; // @[Mux.scala 19:72:@1973.4]
  wire [7:0] _T_4006; // @[Mux.scala 19:72:@1974.4]
  wire [7:0] _T_4013; // @[Mux.scala 19:72:@1981.4]
  wire [7:0] _T_4015; // @[Mux.scala 19:72:@1982.4]
  wire [7:0] _T_4022; // @[Mux.scala 19:72:@1989.4]
  wire [7:0] _T_4024; // @[Mux.scala 19:72:@1990.4]
  wire [7:0] _T_4031; // @[Mux.scala 19:72:@1997.4]
  wire [7:0] _T_4033; // @[Mux.scala 19:72:@1998.4]
  wire [7:0] _T_4040; // @[Mux.scala 19:72:@2005.4]
  wire [7:0] _T_4042; // @[Mux.scala 19:72:@2006.4]
  wire [7:0] _T_4043; // @[Mux.scala 19:72:@2007.4]
  wire [7:0] _T_4044; // @[Mux.scala 19:72:@2008.4]
  wire [7:0] _T_4045; // @[Mux.scala 19:72:@2009.4]
  wire [7:0] _T_4046; // @[Mux.scala 19:72:@2010.4]
  wire [7:0] _T_4047; // @[Mux.scala 19:72:@2011.4]
  wire [7:0] _T_4048; // @[Mux.scala 19:72:@2012.4]
  wire [7:0] _T_4049; // @[Mux.scala 19:72:@2013.4]
  wire  inputAddrPriorityPorts_1_0; // @[Mux.scala 19:72:@2017.4]
  wire  inputAddrPriorityPorts_1_1; // @[Mux.scala 19:72:@2019.4]
  wire  inputAddrPriorityPorts_1_2; // @[Mux.scala 19:72:@2021.4]
  wire  inputAddrPriorityPorts_1_3; // @[Mux.scala 19:72:@2023.4]
  wire  inputAddrPriorityPorts_1_4; // @[Mux.scala 19:72:@2025.4]
  wire  inputAddrPriorityPorts_1_5; // @[Mux.scala 19:72:@2027.4]
  wire  inputAddrPriorityPorts_1_6; // @[Mux.scala 19:72:@2029.4]
  wire  inputAddrPriorityPorts_1_7; // @[Mux.scala 19:72:@2031.4]
  wire [7:0] _T_4163; // @[Mux.scala 31:69:@2061.4]
  wire [7:0] _T_4164; // @[Mux.scala 31:69:@2062.4]
  wire [7:0] _T_4165; // @[Mux.scala 31:69:@2063.4]
  wire [7:0] _T_4166; // @[Mux.scala 31:69:@2064.4]
  wire [7:0] _T_4167; // @[Mux.scala 31:69:@2065.4]
  wire [7:0] _T_4168; // @[Mux.scala 31:69:@2066.4]
  wire [7:0] _T_4169; // @[Mux.scala 31:69:@2067.4]
  wire [7:0] _T_4170; // @[Mux.scala 31:69:@2068.4]
  wire  _T_4171; // @[OneHot.scala 66:30:@2069.4]
  wire  _T_4172; // @[OneHot.scala 66:30:@2070.4]
  wire  _T_4173; // @[OneHot.scala 66:30:@2071.4]
  wire  _T_4174; // @[OneHot.scala 66:30:@2072.4]
  wire  _T_4175; // @[OneHot.scala 66:30:@2073.4]
  wire  _T_4176; // @[OneHot.scala 66:30:@2074.4]
  wire  _T_4177; // @[OneHot.scala 66:30:@2075.4]
  wire  _T_4178; // @[OneHot.scala 66:30:@2076.4]
  wire [7:0] _T_4203; // @[Mux.scala 31:69:@2086.4]
  wire [7:0] _T_4204; // @[Mux.scala 31:69:@2087.4]
  wire [7:0] _T_4205; // @[Mux.scala 31:69:@2088.4]
  wire [7:0] _T_4206; // @[Mux.scala 31:69:@2089.4]
  wire [7:0] _T_4207; // @[Mux.scala 31:69:@2090.4]
  wire [7:0] _T_4208; // @[Mux.scala 31:69:@2091.4]
  wire [7:0] _T_4209; // @[Mux.scala 31:69:@2092.4]
  wire [7:0] _T_4210; // @[Mux.scala 31:69:@2093.4]
  wire  _T_4211; // @[OneHot.scala 66:30:@2094.4]
  wire  _T_4212; // @[OneHot.scala 66:30:@2095.4]
  wire  _T_4213; // @[OneHot.scala 66:30:@2096.4]
  wire  _T_4214; // @[OneHot.scala 66:30:@2097.4]
  wire  _T_4215; // @[OneHot.scala 66:30:@2098.4]
  wire  _T_4216; // @[OneHot.scala 66:30:@2099.4]
  wire  _T_4217; // @[OneHot.scala 66:30:@2100.4]
  wire  _T_4218; // @[OneHot.scala 66:30:@2101.4]
  wire [7:0] _T_4243; // @[Mux.scala 31:69:@2111.4]
  wire [7:0] _T_4244; // @[Mux.scala 31:69:@2112.4]
  wire [7:0] _T_4245; // @[Mux.scala 31:69:@2113.4]
  wire [7:0] _T_4246; // @[Mux.scala 31:69:@2114.4]
  wire [7:0] _T_4247; // @[Mux.scala 31:69:@2115.4]
  wire [7:0] _T_4248; // @[Mux.scala 31:69:@2116.4]
  wire [7:0] _T_4249; // @[Mux.scala 31:69:@2117.4]
  wire [7:0] _T_4250; // @[Mux.scala 31:69:@2118.4]
  wire  _T_4251; // @[OneHot.scala 66:30:@2119.4]
  wire  _T_4252; // @[OneHot.scala 66:30:@2120.4]
  wire  _T_4253; // @[OneHot.scala 66:30:@2121.4]
  wire  _T_4254; // @[OneHot.scala 66:30:@2122.4]
  wire  _T_4255; // @[OneHot.scala 66:30:@2123.4]
  wire  _T_4256; // @[OneHot.scala 66:30:@2124.4]
  wire  _T_4257; // @[OneHot.scala 66:30:@2125.4]
  wire  _T_4258; // @[OneHot.scala 66:30:@2126.4]
  wire [7:0] _T_4283; // @[Mux.scala 31:69:@2136.4]
  wire [7:0] _T_4284; // @[Mux.scala 31:69:@2137.4]
  wire [7:0] _T_4285; // @[Mux.scala 31:69:@2138.4]
  wire [7:0] _T_4286; // @[Mux.scala 31:69:@2139.4]
  wire [7:0] _T_4287; // @[Mux.scala 31:69:@2140.4]
  wire [7:0] _T_4288; // @[Mux.scala 31:69:@2141.4]
  wire [7:0] _T_4289; // @[Mux.scala 31:69:@2142.4]
  wire [7:0] _T_4290; // @[Mux.scala 31:69:@2143.4]
  wire  _T_4291; // @[OneHot.scala 66:30:@2144.4]
  wire  _T_4292; // @[OneHot.scala 66:30:@2145.4]
  wire  _T_4293; // @[OneHot.scala 66:30:@2146.4]
  wire  _T_4294; // @[OneHot.scala 66:30:@2147.4]
  wire  _T_4295; // @[OneHot.scala 66:30:@2148.4]
  wire  _T_4296; // @[OneHot.scala 66:30:@2149.4]
  wire  _T_4297; // @[OneHot.scala 66:30:@2150.4]
  wire  _T_4298; // @[OneHot.scala 66:30:@2151.4]
  wire [7:0] _T_4323; // @[Mux.scala 31:69:@2161.4]
  wire [7:0] _T_4324; // @[Mux.scala 31:69:@2162.4]
  wire [7:0] _T_4325; // @[Mux.scala 31:69:@2163.4]
  wire [7:0] _T_4326; // @[Mux.scala 31:69:@2164.4]
  wire [7:0] _T_4327; // @[Mux.scala 31:69:@2165.4]
  wire [7:0] _T_4328; // @[Mux.scala 31:69:@2166.4]
  wire [7:0] _T_4329; // @[Mux.scala 31:69:@2167.4]
  wire [7:0] _T_4330; // @[Mux.scala 31:69:@2168.4]
  wire  _T_4331; // @[OneHot.scala 66:30:@2169.4]
  wire  _T_4332; // @[OneHot.scala 66:30:@2170.4]
  wire  _T_4333; // @[OneHot.scala 66:30:@2171.4]
  wire  _T_4334; // @[OneHot.scala 66:30:@2172.4]
  wire  _T_4335; // @[OneHot.scala 66:30:@2173.4]
  wire  _T_4336; // @[OneHot.scala 66:30:@2174.4]
  wire  _T_4337; // @[OneHot.scala 66:30:@2175.4]
  wire  _T_4338; // @[OneHot.scala 66:30:@2176.4]
  wire [7:0] _T_4363; // @[Mux.scala 31:69:@2186.4]
  wire [7:0] _T_4364; // @[Mux.scala 31:69:@2187.4]
  wire [7:0] _T_4365; // @[Mux.scala 31:69:@2188.4]
  wire [7:0] _T_4366; // @[Mux.scala 31:69:@2189.4]
  wire [7:0] _T_4367; // @[Mux.scala 31:69:@2190.4]
  wire [7:0] _T_4368; // @[Mux.scala 31:69:@2191.4]
  wire [7:0] _T_4369; // @[Mux.scala 31:69:@2192.4]
  wire [7:0] _T_4370; // @[Mux.scala 31:69:@2193.4]
  wire  _T_4371; // @[OneHot.scala 66:30:@2194.4]
  wire  _T_4372; // @[OneHot.scala 66:30:@2195.4]
  wire  _T_4373; // @[OneHot.scala 66:30:@2196.4]
  wire  _T_4374; // @[OneHot.scala 66:30:@2197.4]
  wire  _T_4375; // @[OneHot.scala 66:30:@2198.4]
  wire  _T_4376; // @[OneHot.scala 66:30:@2199.4]
  wire  _T_4377; // @[OneHot.scala 66:30:@2200.4]
  wire  _T_4378; // @[OneHot.scala 66:30:@2201.4]
  wire [7:0] _T_4403; // @[Mux.scala 31:69:@2211.4]
  wire [7:0] _T_4404; // @[Mux.scala 31:69:@2212.4]
  wire [7:0] _T_4405; // @[Mux.scala 31:69:@2213.4]
  wire [7:0] _T_4406; // @[Mux.scala 31:69:@2214.4]
  wire [7:0] _T_4407; // @[Mux.scala 31:69:@2215.4]
  wire [7:0] _T_4408; // @[Mux.scala 31:69:@2216.4]
  wire [7:0] _T_4409; // @[Mux.scala 31:69:@2217.4]
  wire [7:0] _T_4410; // @[Mux.scala 31:69:@2218.4]
  wire  _T_4411; // @[OneHot.scala 66:30:@2219.4]
  wire  _T_4412; // @[OneHot.scala 66:30:@2220.4]
  wire  _T_4413; // @[OneHot.scala 66:30:@2221.4]
  wire  _T_4414; // @[OneHot.scala 66:30:@2222.4]
  wire  _T_4415; // @[OneHot.scala 66:30:@2223.4]
  wire  _T_4416; // @[OneHot.scala 66:30:@2224.4]
  wire  _T_4417; // @[OneHot.scala 66:30:@2225.4]
  wire  _T_4418; // @[OneHot.scala 66:30:@2226.4]
  wire [7:0] _T_4443; // @[Mux.scala 31:69:@2236.4]
  wire [7:0] _T_4444; // @[Mux.scala 31:69:@2237.4]
  wire [7:0] _T_4445; // @[Mux.scala 31:69:@2238.4]
  wire [7:0] _T_4446; // @[Mux.scala 31:69:@2239.4]
  wire [7:0] _T_4447; // @[Mux.scala 31:69:@2240.4]
  wire [7:0] _T_4448; // @[Mux.scala 31:69:@2241.4]
  wire [7:0] _T_4449; // @[Mux.scala 31:69:@2242.4]
  wire [7:0] _T_4450; // @[Mux.scala 31:69:@2243.4]
  wire  _T_4451; // @[OneHot.scala 66:30:@2244.4]
  wire  _T_4452; // @[OneHot.scala 66:30:@2245.4]
  wire  _T_4453; // @[OneHot.scala 66:30:@2246.4]
  wire  _T_4454; // @[OneHot.scala 66:30:@2247.4]
  wire  _T_4455; // @[OneHot.scala 66:30:@2248.4]
  wire  _T_4456; // @[OneHot.scala 66:30:@2249.4]
  wire  _T_4457; // @[OneHot.scala 66:30:@2250.4]
  wire  _T_4458; // @[OneHot.scala 66:30:@2251.4]
  wire [7:0] _T_4499; // @[Mux.scala 19:72:@2267.4]
  wire [7:0] _T_4501; // @[Mux.scala 19:72:@2268.4]
  wire [7:0] _T_4508; // @[Mux.scala 19:72:@2275.4]
  wire [7:0] _T_4510; // @[Mux.scala 19:72:@2276.4]
  wire [7:0] _T_4517; // @[Mux.scala 19:72:@2283.4]
  wire [7:0] _T_4519; // @[Mux.scala 19:72:@2284.4]
  wire [7:0] _T_4526; // @[Mux.scala 19:72:@2291.4]
  wire [7:0] _T_4528; // @[Mux.scala 19:72:@2292.4]
  wire [7:0] _T_4535; // @[Mux.scala 19:72:@2299.4]
  wire [7:0] _T_4537; // @[Mux.scala 19:72:@2300.4]
  wire [7:0] _T_4544; // @[Mux.scala 19:72:@2307.4]
  wire [7:0] _T_4546; // @[Mux.scala 19:72:@2308.4]
  wire [7:0] _T_4553; // @[Mux.scala 19:72:@2315.4]
  wire [7:0] _T_4555; // @[Mux.scala 19:72:@2316.4]
  wire [7:0] _T_4562; // @[Mux.scala 19:72:@2323.4]
  wire [7:0] _T_4564; // @[Mux.scala 19:72:@2324.4]
  wire [7:0] _T_4565; // @[Mux.scala 19:72:@2325.4]
  wire [7:0] _T_4566; // @[Mux.scala 19:72:@2326.4]
  wire [7:0] _T_4567; // @[Mux.scala 19:72:@2327.4]
  wire [7:0] _T_4568; // @[Mux.scala 19:72:@2328.4]
  wire [7:0] _T_4569; // @[Mux.scala 19:72:@2329.4]
  wire [7:0] _T_4570; // @[Mux.scala 19:72:@2330.4]
  wire [7:0] _T_4571; // @[Mux.scala 19:72:@2331.4]
  wire  inputDataPriorityPorts_1_0; // @[Mux.scala 19:72:@2335.4]
  wire  inputDataPriorityPorts_1_1; // @[Mux.scala 19:72:@2337.4]
  wire  inputDataPriorityPorts_1_2; // @[Mux.scala 19:72:@2339.4]
  wire  inputDataPriorityPorts_1_3; // @[Mux.scala 19:72:@2341.4]
  wire  inputDataPriorityPorts_1_4; // @[Mux.scala 19:72:@2343.4]
  wire  inputDataPriorityPorts_1_5; // @[Mux.scala 19:72:@2345.4]
  wire  inputDataPriorityPorts_1_6; // @[Mux.scala 19:72:@2347.4]
  wire  inputDataPriorityPorts_1_7; // @[Mux.scala 19:72:@2349.4]
  wire  _T_4653; // @[StoreQueue.scala 209:52:@2365.6]
  wire  _T_4654; // @[StoreQueue.scala 209:81:@2366.6]
  wire  _T_4657; // @[StoreQueue.scala 209:52:@2368.6]
  wire  _T_4658; // @[StoreQueue.scala 209:81:@2369.6]
  wire  _T_4669; // @[StoreQueue.scala 210:30:@2374.6]
  wire [1:0] _T_4670; // @[OneHot.scala 18:45:@2376.8]
  wire  _T_4671; // @[CircuitMath.scala 30:8:@2377.8]
  wire [31:0] _GEN_305; // @[StoreQueue.scala 211:30:@2378.8]
  wire [31:0] _GEN_306; // @[StoreQueue.scala 210:40:@2375.6]
  wire  _GEN_307; // @[StoreQueue.scala 210:40:@2375.6]
  wire  _T_4676; // @[StoreQueue.scala 215:52:@2382.6]
  wire  _T_4677; // @[StoreQueue.scala 215:81:@2383.6]
  wire  _T_4680; // @[StoreQueue.scala 215:52:@2385.6]
  wire  _T_4681; // @[StoreQueue.scala 215:81:@2386.6]
  wire  _T_4692; // @[StoreQueue.scala 216:30:@2391.6]
  wire [1:0] _T_4693; // @[OneHot.scala 18:45:@2393.8]
  wire  _T_4694; // @[CircuitMath.scala 30:8:@2394.8]
  wire [31:0] _GEN_309; // @[StoreQueue.scala 217:30:@2395.8]
  wire [31:0] _GEN_310; // @[StoreQueue.scala 216:40:@2392.6]
  wire  _GEN_311; // @[StoreQueue.scala 216:40:@2392.6]
  wire  _GEN_312; // @[StoreQueue.scala 204:35:@2359.4]
  wire  _GEN_313; // @[StoreQueue.scala 204:35:@2359.4]
  wire [31:0] _GEN_314; // @[StoreQueue.scala 204:35:@2359.4]
  wire [31:0] _GEN_315; // @[StoreQueue.scala 204:35:@2359.4]
  wire  _T_4701; // @[StoreQueue.scala 209:52:@2405.6]
  wire  _T_4702; // @[StoreQueue.scala 209:81:@2406.6]
  wire  _T_4705; // @[StoreQueue.scala 209:52:@2408.6]
  wire  _T_4706; // @[StoreQueue.scala 209:81:@2409.6]
  wire  _T_4717; // @[StoreQueue.scala 210:30:@2414.6]
  wire [1:0] _T_4718; // @[OneHot.scala 18:45:@2416.8]
  wire  _T_4719; // @[CircuitMath.scala 30:8:@2417.8]
  wire [31:0] _GEN_317; // @[StoreQueue.scala 211:30:@2418.8]
  wire [31:0] _GEN_318; // @[StoreQueue.scala 210:40:@2415.6]
  wire  _GEN_319; // @[StoreQueue.scala 210:40:@2415.6]
  wire  _T_4724; // @[StoreQueue.scala 215:52:@2422.6]
  wire  _T_4725; // @[StoreQueue.scala 215:81:@2423.6]
  wire  _T_4728; // @[StoreQueue.scala 215:52:@2425.6]
  wire  _T_4729; // @[StoreQueue.scala 215:81:@2426.6]
  wire  _T_4740; // @[StoreQueue.scala 216:30:@2431.6]
  wire [1:0] _T_4741; // @[OneHot.scala 18:45:@2433.8]
  wire  _T_4742; // @[CircuitMath.scala 30:8:@2434.8]
  wire [31:0] _GEN_321; // @[StoreQueue.scala 217:30:@2435.8]
  wire [31:0] _GEN_322; // @[StoreQueue.scala 216:40:@2432.6]
  wire  _GEN_323; // @[StoreQueue.scala 216:40:@2432.6]
  wire  _GEN_324; // @[StoreQueue.scala 204:35:@2399.4]
  wire  _GEN_325; // @[StoreQueue.scala 204:35:@2399.4]
  wire [31:0] _GEN_326; // @[StoreQueue.scala 204:35:@2399.4]
  wire [31:0] _GEN_327; // @[StoreQueue.scala 204:35:@2399.4]
  wire  _T_4749; // @[StoreQueue.scala 209:52:@2445.6]
  wire  _T_4750; // @[StoreQueue.scala 209:81:@2446.6]
  wire  _T_4753; // @[StoreQueue.scala 209:52:@2448.6]
  wire  _T_4754; // @[StoreQueue.scala 209:81:@2449.6]
  wire  _T_4765; // @[StoreQueue.scala 210:30:@2454.6]
  wire [1:0] _T_4766; // @[OneHot.scala 18:45:@2456.8]
  wire  _T_4767; // @[CircuitMath.scala 30:8:@2457.8]
  wire [31:0] _GEN_329; // @[StoreQueue.scala 211:30:@2458.8]
  wire [31:0] _GEN_330; // @[StoreQueue.scala 210:40:@2455.6]
  wire  _GEN_331; // @[StoreQueue.scala 210:40:@2455.6]
  wire  _T_4772; // @[StoreQueue.scala 215:52:@2462.6]
  wire  _T_4773; // @[StoreQueue.scala 215:81:@2463.6]
  wire  _T_4776; // @[StoreQueue.scala 215:52:@2465.6]
  wire  _T_4777; // @[StoreQueue.scala 215:81:@2466.6]
  wire  _T_4788; // @[StoreQueue.scala 216:30:@2471.6]
  wire [1:0] _T_4789; // @[OneHot.scala 18:45:@2473.8]
  wire  _T_4790; // @[CircuitMath.scala 30:8:@2474.8]
  wire [31:0] _GEN_333; // @[StoreQueue.scala 217:30:@2475.8]
  wire [31:0] _GEN_334; // @[StoreQueue.scala 216:40:@2472.6]
  wire  _GEN_335; // @[StoreQueue.scala 216:40:@2472.6]
  wire  _GEN_336; // @[StoreQueue.scala 204:35:@2439.4]
  wire  _GEN_337; // @[StoreQueue.scala 204:35:@2439.4]
  wire [31:0] _GEN_338; // @[StoreQueue.scala 204:35:@2439.4]
  wire [31:0] _GEN_339; // @[StoreQueue.scala 204:35:@2439.4]
  wire  _T_4797; // @[StoreQueue.scala 209:52:@2485.6]
  wire  _T_4798; // @[StoreQueue.scala 209:81:@2486.6]
  wire  _T_4801; // @[StoreQueue.scala 209:52:@2488.6]
  wire  _T_4802; // @[StoreQueue.scala 209:81:@2489.6]
  wire  _T_4813; // @[StoreQueue.scala 210:30:@2494.6]
  wire [1:0] _T_4814; // @[OneHot.scala 18:45:@2496.8]
  wire  _T_4815; // @[CircuitMath.scala 30:8:@2497.8]
  wire [31:0] _GEN_341; // @[StoreQueue.scala 211:30:@2498.8]
  wire [31:0] _GEN_342; // @[StoreQueue.scala 210:40:@2495.6]
  wire  _GEN_343; // @[StoreQueue.scala 210:40:@2495.6]
  wire  _T_4820; // @[StoreQueue.scala 215:52:@2502.6]
  wire  _T_4821; // @[StoreQueue.scala 215:81:@2503.6]
  wire  _T_4824; // @[StoreQueue.scala 215:52:@2505.6]
  wire  _T_4825; // @[StoreQueue.scala 215:81:@2506.6]
  wire  _T_4836; // @[StoreQueue.scala 216:30:@2511.6]
  wire [1:0] _T_4837; // @[OneHot.scala 18:45:@2513.8]
  wire  _T_4838; // @[CircuitMath.scala 30:8:@2514.8]
  wire [31:0] _GEN_345; // @[StoreQueue.scala 217:30:@2515.8]
  wire [31:0] _GEN_346; // @[StoreQueue.scala 216:40:@2512.6]
  wire  _GEN_347; // @[StoreQueue.scala 216:40:@2512.6]
  wire  _GEN_348; // @[StoreQueue.scala 204:35:@2479.4]
  wire  _GEN_349; // @[StoreQueue.scala 204:35:@2479.4]
  wire [31:0] _GEN_350; // @[StoreQueue.scala 204:35:@2479.4]
  wire [31:0] _GEN_351; // @[StoreQueue.scala 204:35:@2479.4]
  wire  _T_4845; // @[StoreQueue.scala 209:52:@2525.6]
  wire  _T_4846; // @[StoreQueue.scala 209:81:@2526.6]
  wire  _T_4849; // @[StoreQueue.scala 209:52:@2528.6]
  wire  _T_4850; // @[StoreQueue.scala 209:81:@2529.6]
  wire  _T_4861; // @[StoreQueue.scala 210:30:@2534.6]
  wire [1:0] _T_4862; // @[OneHot.scala 18:45:@2536.8]
  wire  _T_4863; // @[CircuitMath.scala 30:8:@2537.8]
  wire [31:0] _GEN_353; // @[StoreQueue.scala 211:30:@2538.8]
  wire [31:0] _GEN_354; // @[StoreQueue.scala 210:40:@2535.6]
  wire  _GEN_355; // @[StoreQueue.scala 210:40:@2535.6]
  wire  _T_4868; // @[StoreQueue.scala 215:52:@2542.6]
  wire  _T_4869; // @[StoreQueue.scala 215:81:@2543.6]
  wire  _T_4872; // @[StoreQueue.scala 215:52:@2545.6]
  wire  _T_4873; // @[StoreQueue.scala 215:81:@2546.6]
  wire  _T_4884; // @[StoreQueue.scala 216:30:@2551.6]
  wire [1:0] _T_4885; // @[OneHot.scala 18:45:@2553.8]
  wire  _T_4886; // @[CircuitMath.scala 30:8:@2554.8]
  wire [31:0] _GEN_357; // @[StoreQueue.scala 217:30:@2555.8]
  wire [31:0] _GEN_358; // @[StoreQueue.scala 216:40:@2552.6]
  wire  _GEN_359; // @[StoreQueue.scala 216:40:@2552.6]
  wire  _GEN_360; // @[StoreQueue.scala 204:35:@2519.4]
  wire  _GEN_361; // @[StoreQueue.scala 204:35:@2519.4]
  wire [31:0] _GEN_362; // @[StoreQueue.scala 204:35:@2519.4]
  wire [31:0] _GEN_363; // @[StoreQueue.scala 204:35:@2519.4]
  wire  _T_4893; // @[StoreQueue.scala 209:52:@2565.6]
  wire  _T_4894; // @[StoreQueue.scala 209:81:@2566.6]
  wire  _T_4897; // @[StoreQueue.scala 209:52:@2568.6]
  wire  _T_4898; // @[StoreQueue.scala 209:81:@2569.6]
  wire  _T_4909; // @[StoreQueue.scala 210:30:@2574.6]
  wire [1:0] _T_4910; // @[OneHot.scala 18:45:@2576.8]
  wire  _T_4911; // @[CircuitMath.scala 30:8:@2577.8]
  wire [31:0] _GEN_365; // @[StoreQueue.scala 211:30:@2578.8]
  wire [31:0] _GEN_366; // @[StoreQueue.scala 210:40:@2575.6]
  wire  _GEN_367; // @[StoreQueue.scala 210:40:@2575.6]
  wire  _T_4916; // @[StoreQueue.scala 215:52:@2582.6]
  wire  _T_4917; // @[StoreQueue.scala 215:81:@2583.6]
  wire  _T_4920; // @[StoreQueue.scala 215:52:@2585.6]
  wire  _T_4921; // @[StoreQueue.scala 215:81:@2586.6]
  wire  _T_4932; // @[StoreQueue.scala 216:30:@2591.6]
  wire [1:0] _T_4933; // @[OneHot.scala 18:45:@2593.8]
  wire  _T_4934; // @[CircuitMath.scala 30:8:@2594.8]
  wire [31:0] _GEN_369; // @[StoreQueue.scala 217:30:@2595.8]
  wire [31:0] _GEN_370; // @[StoreQueue.scala 216:40:@2592.6]
  wire  _GEN_371; // @[StoreQueue.scala 216:40:@2592.6]
  wire  _GEN_372; // @[StoreQueue.scala 204:35:@2559.4]
  wire  _GEN_373; // @[StoreQueue.scala 204:35:@2559.4]
  wire [31:0] _GEN_374; // @[StoreQueue.scala 204:35:@2559.4]
  wire [31:0] _GEN_375; // @[StoreQueue.scala 204:35:@2559.4]
  wire  _T_4941; // @[StoreQueue.scala 209:52:@2605.6]
  wire  _T_4942; // @[StoreQueue.scala 209:81:@2606.6]
  wire  _T_4945; // @[StoreQueue.scala 209:52:@2608.6]
  wire  _T_4946; // @[StoreQueue.scala 209:81:@2609.6]
  wire  _T_4957; // @[StoreQueue.scala 210:30:@2614.6]
  wire [1:0] _T_4958; // @[OneHot.scala 18:45:@2616.8]
  wire  _T_4959; // @[CircuitMath.scala 30:8:@2617.8]
  wire [31:0] _GEN_377; // @[StoreQueue.scala 211:30:@2618.8]
  wire [31:0] _GEN_378; // @[StoreQueue.scala 210:40:@2615.6]
  wire  _GEN_379; // @[StoreQueue.scala 210:40:@2615.6]
  wire  _T_4964; // @[StoreQueue.scala 215:52:@2622.6]
  wire  _T_4965; // @[StoreQueue.scala 215:81:@2623.6]
  wire  _T_4968; // @[StoreQueue.scala 215:52:@2625.6]
  wire  _T_4969; // @[StoreQueue.scala 215:81:@2626.6]
  wire  _T_4980; // @[StoreQueue.scala 216:30:@2631.6]
  wire [1:0] _T_4981; // @[OneHot.scala 18:45:@2633.8]
  wire  _T_4982; // @[CircuitMath.scala 30:8:@2634.8]
  wire [31:0] _GEN_381; // @[StoreQueue.scala 217:30:@2635.8]
  wire [31:0] _GEN_382; // @[StoreQueue.scala 216:40:@2632.6]
  wire  _GEN_383; // @[StoreQueue.scala 216:40:@2632.6]
  wire  _GEN_384; // @[StoreQueue.scala 204:35:@2599.4]
  wire  _GEN_385; // @[StoreQueue.scala 204:35:@2599.4]
  wire [31:0] _GEN_386; // @[StoreQueue.scala 204:35:@2599.4]
  wire [31:0] _GEN_387; // @[StoreQueue.scala 204:35:@2599.4]
  wire  _T_4989; // @[StoreQueue.scala 209:52:@2645.6]
  wire  _T_4990; // @[StoreQueue.scala 209:81:@2646.6]
  wire  _T_4993; // @[StoreQueue.scala 209:52:@2648.6]
  wire  _T_4994; // @[StoreQueue.scala 209:81:@2649.6]
  wire  _T_5005; // @[StoreQueue.scala 210:30:@2654.6]
  wire [1:0] _T_5006; // @[OneHot.scala 18:45:@2656.8]
  wire  _T_5007; // @[CircuitMath.scala 30:8:@2657.8]
  wire [31:0] _GEN_389; // @[StoreQueue.scala 211:30:@2658.8]
  wire [31:0] _GEN_390; // @[StoreQueue.scala 210:40:@2655.6]
  wire  _GEN_391; // @[StoreQueue.scala 210:40:@2655.6]
  wire  _T_5012; // @[StoreQueue.scala 215:52:@2662.6]
  wire  _T_5013; // @[StoreQueue.scala 215:81:@2663.6]
  wire  _T_5016; // @[StoreQueue.scala 215:52:@2665.6]
  wire  _T_5017; // @[StoreQueue.scala 215:81:@2666.6]
  wire  _T_5028; // @[StoreQueue.scala 216:30:@2671.6]
  wire [1:0] _T_5029; // @[OneHot.scala 18:45:@2673.8]
  wire  _T_5030; // @[CircuitMath.scala 30:8:@2674.8]
  wire [31:0] _GEN_393; // @[StoreQueue.scala 217:30:@2675.8]
  wire [31:0] _GEN_394; // @[StoreQueue.scala 216:40:@2672.6]
  wire  _GEN_395; // @[StoreQueue.scala 216:40:@2672.6]
  wire  _GEN_396; // @[StoreQueue.scala 204:35:@2639.4]
  wire  _GEN_397; // @[StoreQueue.scala 204:35:@2639.4]
  wire [31:0] _GEN_398; // @[StoreQueue.scala 204:35:@2639.4]
  wire [31:0] _GEN_399; // @[StoreQueue.scala 204:35:@2639.4]
  wire  _T_5033; // @[StoreQueue.scala 229:23:@2679.4]
  wire [3:0] _T_5036; // @[util.scala 10:8:@2681.6]
  wire [3:0] _GEN_144; // @[util.scala 10:14:@2682.6]
  wire [3:0] _T_5037; // @[util.scala 10:14:@2682.6]
  wire [3:0] _GEN_400; // @[StoreQueue.scala 229:50:@2680.4]
  wire [2:0] _GEN_458; // @[util.scala 10:8:@2686.6]
  wire [3:0] _T_5039; // @[util.scala 10:8:@2686.6]
  wire [3:0] _GEN_145; // @[util.scala 10:14:@2687.6]
  wire [3:0] _T_5040; // @[util.scala 10:14:@2687.6]
  wire [3:0] _GEN_401; // @[StoreQueue.scala 233:20:@2685.4]
  wire  _T_5042; // @[StoreQueue.scala 237:84:@2690.4]
  wire  _T_5043; // @[StoreQueue.scala 237:81:@2691.4]
  wire  _T_5045; // @[StoreQueue.scala 237:84:@2692.4]
  wire  _T_5046; // @[StoreQueue.scala 237:81:@2693.4]
  wire  _T_5048; // @[StoreQueue.scala 237:84:@2694.4]
  wire  _T_5049; // @[StoreQueue.scala 237:81:@2695.4]
  wire  _T_5051; // @[StoreQueue.scala 237:84:@2696.4]
  wire  _T_5052; // @[StoreQueue.scala 237:81:@2697.4]
  wire  _T_5054; // @[StoreQueue.scala 237:84:@2698.4]
  wire  _T_5055; // @[StoreQueue.scala 237:81:@2699.4]
  wire  _T_5057; // @[StoreQueue.scala 237:84:@2700.4]
  wire  _T_5058; // @[StoreQueue.scala 237:81:@2701.4]
  wire  _T_5060; // @[StoreQueue.scala 237:84:@2702.4]
  wire  _T_5061; // @[StoreQueue.scala 237:81:@2703.4]
  wire  _T_5063; // @[StoreQueue.scala 237:84:@2704.4]
  wire  _T_5064; // @[StoreQueue.scala 237:81:@2705.4]
  wire  _T_5081; // @[StoreQueue.scala 237:98:@2716.4]
  wire  _T_5082; // @[StoreQueue.scala 237:98:@2717.4]
  wire  _T_5083; // @[StoreQueue.scala 237:98:@2718.4]
  wire  _T_5084; // @[StoreQueue.scala 237:98:@2719.4]
  wire  _T_5085; // @[StoreQueue.scala 237:98:@2720.4]
  wire  _T_5086; // @[StoreQueue.scala 237:98:@2721.4]
  wire [31:0] _GEN_403; // @[StoreQueue.scala 252:21:@2759.4]
  wire [31:0] _GEN_404; // @[StoreQueue.scala 252:21:@2759.4]
  wire [31:0] _GEN_405; // @[StoreQueue.scala 252:21:@2759.4]
  wire [31:0] _GEN_406; // @[StoreQueue.scala 252:21:@2759.4]
  wire [31:0] _GEN_407; // @[StoreQueue.scala 252:21:@2759.4]
  wire [31:0] _GEN_408; // @[StoreQueue.scala 252:21:@2759.4]
  assign _GEN_410 = {{2'd0}, tail}; // @[util.scala 14:20:@101.4]
  assign _T_956 = 5'h8 - _GEN_410; // @[util.scala 14:20:@101.4]
  assign _T_957 = $unsigned(_T_956); // @[util.scala 14:20:@102.4]
  assign _T_958 = _T_957[4:0]; // @[util.scala 14:20:@103.4]
  assign _GEN_0 = _T_958 % 5'h8; // @[util.scala 14:25:@104.4]
  assign _T_959 = _GEN_0[3:0]; // @[util.scala 14:25:@104.4]
  assign _GEN_411 = {{2'd0}, io_bbNumStores}; // @[StoreQueue.scala 70:46:@105.4]
  assign _T_960 = _T_959 < _GEN_411; // @[StoreQueue.scala 70:46:@105.4]
  assign initBits_0 = _T_960 & io_bbStart; // @[StoreQueue.scala 70:64:@106.4]
  assign _T_965 = 5'h9 - _GEN_410; // @[util.scala 14:20:@108.4]
  assign _T_966 = $unsigned(_T_965); // @[util.scala 14:20:@109.4]
  assign _T_967 = _T_966[4:0]; // @[util.scala 14:20:@110.4]
  assign _GEN_8 = _T_967 % 5'h8; // @[util.scala 14:25:@111.4]
  assign _T_968 = _GEN_8[3:0]; // @[util.scala 14:25:@111.4]
  assign _T_969 = _T_968 < _GEN_411; // @[StoreQueue.scala 70:46:@112.4]
  assign initBits_1 = _T_969 & io_bbStart; // @[StoreQueue.scala 70:64:@113.4]
  assign _T_974 = 5'ha - _GEN_410; // @[util.scala 14:20:@115.4]
  assign _T_975 = $unsigned(_T_974); // @[util.scala 14:20:@116.4]
  assign _T_976 = _T_975[4:0]; // @[util.scala 14:20:@117.4]
  assign _GEN_18 = _T_976 % 5'h8; // @[util.scala 14:25:@118.4]
  assign _T_977 = _GEN_18[3:0]; // @[util.scala 14:25:@118.4]
  assign _T_978 = _T_977 < _GEN_411; // @[StoreQueue.scala 70:46:@119.4]
  assign initBits_2 = _T_978 & io_bbStart; // @[StoreQueue.scala 70:64:@120.4]
  assign _T_983 = 5'hb - _GEN_410; // @[util.scala 14:20:@122.4]
  assign _T_984 = $unsigned(_T_983); // @[util.scala 14:20:@123.4]
  assign _T_985 = _T_984[4:0]; // @[util.scala 14:20:@124.4]
  assign _GEN_26 = _T_985 % 5'h8; // @[util.scala 14:25:@125.4]
  assign _T_986 = _GEN_26[3:0]; // @[util.scala 14:25:@125.4]
  assign _T_987 = _T_986 < _GEN_411; // @[StoreQueue.scala 70:46:@126.4]
  assign initBits_3 = _T_987 & io_bbStart; // @[StoreQueue.scala 70:64:@127.4]
  assign _T_992 = 5'hc - _GEN_410; // @[util.scala 14:20:@129.4]
  assign _T_993 = $unsigned(_T_992); // @[util.scala 14:20:@130.4]
  assign _T_994 = _T_993[4:0]; // @[util.scala 14:20:@131.4]
  assign _GEN_36 = _T_994 % 5'h8; // @[util.scala 14:25:@132.4]
  assign _T_995 = _GEN_36[3:0]; // @[util.scala 14:25:@132.4]
  assign _T_996 = _T_995 < _GEN_411; // @[StoreQueue.scala 70:46:@133.4]
  assign initBits_4 = _T_996 & io_bbStart; // @[StoreQueue.scala 70:64:@134.4]
  assign _T_1001 = 5'hd - _GEN_410; // @[util.scala 14:20:@136.4]
  assign _T_1002 = $unsigned(_T_1001); // @[util.scala 14:20:@137.4]
  assign _T_1003 = _T_1002[4:0]; // @[util.scala 14:20:@138.4]
  assign _GEN_44 = _T_1003 % 5'h8; // @[util.scala 14:25:@139.4]
  assign _T_1004 = _GEN_44[3:0]; // @[util.scala 14:25:@139.4]
  assign _T_1005 = _T_1004 < _GEN_411; // @[StoreQueue.scala 70:46:@140.4]
  assign initBits_5 = _T_1005 & io_bbStart; // @[StoreQueue.scala 70:64:@141.4]
  assign _T_1010 = 5'he - _GEN_410; // @[util.scala 14:20:@143.4]
  assign _T_1011 = $unsigned(_T_1010); // @[util.scala 14:20:@144.4]
  assign _T_1012 = _T_1011[4:0]; // @[util.scala 14:20:@145.4]
  assign _GEN_54 = _T_1012 % 5'h8; // @[util.scala 14:25:@146.4]
  assign _T_1013 = _GEN_54[3:0]; // @[util.scala 14:25:@146.4]
  assign _T_1014 = _T_1013 < _GEN_411; // @[StoreQueue.scala 70:46:@147.4]
  assign initBits_6 = _T_1014 & io_bbStart; // @[StoreQueue.scala 70:64:@148.4]
  assign _T_1019 = 5'hf - _GEN_410; // @[util.scala 14:20:@150.4]
  assign _T_1020 = $unsigned(_T_1019); // @[util.scala 14:20:@151.4]
  assign _T_1021 = _T_1020[4:0]; // @[util.scala 14:20:@152.4]
  assign _GEN_62 = _T_1021 % 5'h8; // @[util.scala 14:25:@153.4]
  assign _T_1022 = _GEN_62[3:0]; // @[util.scala 14:25:@153.4]
  assign _T_1023 = _T_1022 < _GEN_411; // @[StoreQueue.scala 70:46:@154.4]
  assign initBits_7 = _T_1023 & io_bbStart; // @[StoreQueue.scala 70:64:@155.4]
  assign _T_1038 = allocatedEntries_0 | initBits_0; // @[StoreQueue.scala 72:78:@165.4]
  assign _T_1039 = allocatedEntries_1 | initBits_1; // @[StoreQueue.scala 72:78:@166.4]
  assign _T_1040 = allocatedEntries_2 | initBits_2; // @[StoreQueue.scala 72:78:@167.4]
  assign _T_1041 = allocatedEntries_3 | initBits_3; // @[StoreQueue.scala 72:78:@168.4]
  assign _T_1042 = allocatedEntries_4 | initBits_4; // @[StoreQueue.scala 72:78:@169.4]
  assign _T_1043 = allocatedEntries_5 | initBits_5; // @[StoreQueue.scala 72:78:@170.4]
  assign _T_1044 = allocatedEntries_6 | initBits_6; // @[StoreQueue.scala 72:78:@171.4]
  assign _T_1045 = allocatedEntries_7 | initBits_7; // @[StoreQueue.scala 72:78:@172.4]
  assign _T_1068 = _T_959[2:0]; // @[:@196.6]
  assign _GEN_1 = 3'h1 == _T_1068 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_2 = 3'h2 == _T_1068 ? io_bbStoreOffsets_2 : _GEN_1; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_3 = 3'h3 == _T_1068 ? io_bbStoreOffsets_3 : _GEN_2; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_4 = 3'h4 == _T_1068 ? io_bbStoreOffsets_4 : _GEN_3; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_5 = 3'h5 == _T_1068 ? io_bbStoreOffsets_5 : _GEN_4; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_6 = 3'h6 == _T_1068 ? io_bbStoreOffsets_6 : _GEN_5; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_7 = 3'h7 == _T_1068 ? io_bbStoreOffsets_7 : _GEN_6; // @[StoreQueue.scala 76:20:@197.6]
  assign _GEN_9 = 3'h1 == _T_1068 ? io_bbStorePorts_1 : 1'h0; // @[StoreQueue.scala 77:18:@204.6]
  assign _GEN_10 = 3'h2 == _T_1068 ? 1'h0 : _GEN_9; // @[StoreQueue.scala 77:18:@204.6]
  assign _GEN_11 = 3'h3 == _T_1068 ? 1'h0 : _GEN_10; // @[StoreQueue.scala 77:18:@204.6]
  assign _GEN_12 = 3'h4 == _T_1068 ? 1'h0 : _GEN_11; // @[StoreQueue.scala 77:18:@204.6]
  assign _GEN_13 = 3'h5 == _T_1068 ? 1'h0 : _GEN_12; // @[StoreQueue.scala 77:18:@204.6]
  assign _GEN_14 = 3'h6 == _T_1068 ? 1'h0 : _GEN_13; // @[StoreQueue.scala 77:18:@204.6]
  assign _GEN_15 = 3'h7 == _T_1068 ? 1'h0 : _GEN_14; // @[StoreQueue.scala 77:18:@204.6]
  assign _GEN_16 = initBits_0 ? _GEN_7 : offsetQ_0; // @[StoreQueue.scala 75:25:@190.4]
  assign _GEN_17 = initBits_0 ? _GEN_15 : portQ_0; // @[StoreQueue.scala 75:25:@190.4]
  assign _T_1086 = _T_968[2:0]; // @[:@212.6]
  assign _GEN_19 = 3'h1 == _T_1086 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_20 = 3'h2 == _T_1086 ? io_bbStoreOffsets_2 : _GEN_19; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_21 = 3'h3 == _T_1086 ? io_bbStoreOffsets_3 : _GEN_20; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_22 = 3'h4 == _T_1086 ? io_bbStoreOffsets_4 : _GEN_21; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_23 = 3'h5 == _T_1086 ? io_bbStoreOffsets_5 : _GEN_22; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_24 = 3'h6 == _T_1086 ? io_bbStoreOffsets_6 : _GEN_23; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_25 = 3'h7 == _T_1086 ? io_bbStoreOffsets_7 : _GEN_24; // @[StoreQueue.scala 76:20:@213.6]
  assign _GEN_27 = 3'h1 == _T_1086 ? io_bbStorePorts_1 : 1'h0; // @[StoreQueue.scala 77:18:@220.6]
  assign _GEN_28 = 3'h2 == _T_1086 ? 1'h0 : _GEN_27; // @[StoreQueue.scala 77:18:@220.6]
  assign _GEN_29 = 3'h3 == _T_1086 ? 1'h0 : _GEN_28; // @[StoreQueue.scala 77:18:@220.6]
  assign _GEN_30 = 3'h4 == _T_1086 ? 1'h0 : _GEN_29; // @[StoreQueue.scala 77:18:@220.6]
  assign _GEN_31 = 3'h5 == _T_1086 ? 1'h0 : _GEN_30; // @[StoreQueue.scala 77:18:@220.6]
  assign _GEN_32 = 3'h6 == _T_1086 ? 1'h0 : _GEN_31; // @[StoreQueue.scala 77:18:@220.6]
  assign _GEN_33 = 3'h7 == _T_1086 ? 1'h0 : _GEN_32; // @[StoreQueue.scala 77:18:@220.6]
  assign _GEN_34 = initBits_1 ? _GEN_25 : offsetQ_1; // @[StoreQueue.scala 75:25:@206.4]
  assign _GEN_35 = initBits_1 ? _GEN_33 : portQ_1; // @[StoreQueue.scala 75:25:@206.4]
  assign _T_1104 = _T_977[2:0]; // @[:@228.6]
  assign _GEN_37 = 3'h1 == _T_1104 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_38 = 3'h2 == _T_1104 ? io_bbStoreOffsets_2 : _GEN_37; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_39 = 3'h3 == _T_1104 ? io_bbStoreOffsets_3 : _GEN_38; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_40 = 3'h4 == _T_1104 ? io_bbStoreOffsets_4 : _GEN_39; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_41 = 3'h5 == _T_1104 ? io_bbStoreOffsets_5 : _GEN_40; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_42 = 3'h6 == _T_1104 ? io_bbStoreOffsets_6 : _GEN_41; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_43 = 3'h7 == _T_1104 ? io_bbStoreOffsets_7 : _GEN_42; // @[StoreQueue.scala 76:20:@229.6]
  assign _GEN_45 = 3'h1 == _T_1104 ? io_bbStorePorts_1 : 1'h0; // @[StoreQueue.scala 77:18:@236.6]
  assign _GEN_46 = 3'h2 == _T_1104 ? 1'h0 : _GEN_45; // @[StoreQueue.scala 77:18:@236.6]
  assign _GEN_47 = 3'h3 == _T_1104 ? 1'h0 : _GEN_46; // @[StoreQueue.scala 77:18:@236.6]
  assign _GEN_48 = 3'h4 == _T_1104 ? 1'h0 : _GEN_47; // @[StoreQueue.scala 77:18:@236.6]
  assign _GEN_49 = 3'h5 == _T_1104 ? 1'h0 : _GEN_48; // @[StoreQueue.scala 77:18:@236.6]
  assign _GEN_50 = 3'h6 == _T_1104 ? 1'h0 : _GEN_49; // @[StoreQueue.scala 77:18:@236.6]
  assign _GEN_51 = 3'h7 == _T_1104 ? 1'h0 : _GEN_50; // @[StoreQueue.scala 77:18:@236.6]
  assign _GEN_52 = initBits_2 ? _GEN_43 : offsetQ_2; // @[StoreQueue.scala 75:25:@222.4]
  assign _GEN_53 = initBits_2 ? _GEN_51 : portQ_2; // @[StoreQueue.scala 75:25:@222.4]
  assign _T_1122 = _T_986[2:0]; // @[:@244.6]
  assign _GEN_55 = 3'h1 == _T_1122 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_56 = 3'h2 == _T_1122 ? io_bbStoreOffsets_2 : _GEN_55; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_57 = 3'h3 == _T_1122 ? io_bbStoreOffsets_3 : _GEN_56; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_58 = 3'h4 == _T_1122 ? io_bbStoreOffsets_4 : _GEN_57; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_59 = 3'h5 == _T_1122 ? io_bbStoreOffsets_5 : _GEN_58; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_60 = 3'h6 == _T_1122 ? io_bbStoreOffsets_6 : _GEN_59; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_61 = 3'h7 == _T_1122 ? io_bbStoreOffsets_7 : _GEN_60; // @[StoreQueue.scala 76:20:@245.6]
  assign _GEN_63 = 3'h1 == _T_1122 ? io_bbStorePorts_1 : 1'h0; // @[StoreQueue.scala 77:18:@252.6]
  assign _GEN_64 = 3'h2 == _T_1122 ? 1'h0 : _GEN_63; // @[StoreQueue.scala 77:18:@252.6]
  assign _GEN_65 = 3'h3 == _T_1122 ? 1'h0 : _GEN_64; // @[StoreQueue.scala 77:18:@252.6]
  assign _GEN_66 = 3'h4 == _T_1122 ? 1'h0 : _GEN_65; // @[StoreQueue.scala 77:18:@252.6]
  assign _GEN_67 = 3'h5 == _T_1122 ? 1'h0 : _GEN_66; // @[StoreQueue.scala 77:18:@252.6]
  assign _GEN_68 = 3'h6 == _T_1122 ? 1'h0 : _GEN_67; // @[StoreQueue.scala 77:18:@252.6]
  assign _GEN_69 = 3'h7 == _T_1122 ? 1'h0 : _GEN_68; // @[StoreQueue.scala 77:18:@252.6]
  assign _GEN_70 = initBits_3 ? _GEN_61 : offsetQ_3; // @[StoreQueue.scala 75:25:@238.4]
  assign _GEN_71 = initBits_3 ? _GEN_69 : portQ_3; // @[StoreQueue.scala 75:25:@238.4]
  assign _T_1140 = _T_995[2:0]; // @[:@260.6]
  assign _GEN_73 = 3'h1 == _T_1140 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_74 = 3'h2 == _T_1140 ? io_bbStoreOffsets_2 : _GEN_73; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_75 = 3'h3 == _T_1140 ? io_bbStoreOffsets_3 : _GEN_74; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_76 = 3'h4 == _T_1140 ? io_bbStoreOffsets_4 : _GEN_75; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_77 = 3'h5 == _T_1140 ? io_bbStoreOffsets_5 : _GEN_76; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_78 = 3'h6 == _T_1140 ? io_bbStoreOffsets_6 : _GEN_77; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_79 = 3'h7 == _T_1140 ? io_bbStoreOffsets_7 : _GEN_78; // @[StoreQueue.scala 76:20:@261.6]
  assign _GEN_81 = 3'h1 == _T_1140 ? io_bbStorePorts_1 : 1'h0; // @[StoreQueue.scala 77:18:@268.6]
  assign _GEN_82 = 3'h2 == _T_1140 ? 1'h0 : _GEN_81; // @[StoreQueue.scala 77:18:@268.6]
  assign _GEN_83 = 3'h3 == _T_1140 ? 1'h0 : _GEN_82; // @[StoreQueue.scala 77:18:@268.6]
  assign _GEN_84 = 3'h4 == _T_1140 ? 1'h0 : _GEN_83; // @[StoreQueue.scala 77:18:@268.6]
  assign _GEN_85 = 3'h5 == _T_1140 ? 1'h0 : _GEN_84; // @[StoreQueue.scala 77:18:@268.6]
  assign _GEN_86 = 3'h6 == _T_1140 ? 1'h0 : _GEN_85; // @[StoreQueue.scala 77:18:@268.6]
  assign _GEN_87 = 3'h7 == _T_1140 ? 1'h0 : _GEN_86; // @[StoreQueue.scala 77:18:@268.6]
  assign _GEN_88 = initBits_4 ? _GEN_79 : offsetQ_4; // @[StoreQueue.scala 75:25:@254.4]
  assign _GEN_89 = initBits_4 ? _GEN_87 : portQ_4; // @[StoreQueue.scala 75:25:@254.4]
  assign _T_1158 = _T_1004[2:0]; // @[:@276.6]
  assign _GEN_91 = 3'h1 == _T_1158 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_92 = 3'h2 == _T_1158 ? io_bbStoreOffsets_2 : _GEN_91; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_93 = 3'h3 == _T_1158 ? io_bbStoreOffsets_3 : _GEN_92; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_94 = 3'h4 == _T_1158 ? io_bbStoreOffsets_4 : _GEN_93; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_95 = 3'h5 == _T_1158 ? io_bbStoreOffsets_5 : _GEN_94; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_96 = 3'h6 == _T_1158 ? io_bbStoreOffsets_6 : _GEN_95; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_97 = 3'h7 == _T_1158 ? io_bbStoreOffsets_7 : _GEN_96; // @[StoreQueue.scala 76:20:@277.6]
  assign _GEN_99 = 3'h1 == _T_1158 ? io_bbStorePorts_1 : 1'h0; // @[StoreQueue.scala 77:18:@284.6]
  assign _GEN_100 = 3'h2 == _T_1158 ? 1'h0 : _GEN_99; // @[StoreQueue.scala 77:18:@284.6]
  assign _GEN_101 = 3'h3 == _T_1158 ? 1'h0 : _GEN_100; // @[StoreQueue.scala 77:18:@284.6]
  assign _GEN_102 = 3'h4 == _T_1158 ? 1'h0 : _GEN_101; // @[StoreQueue.scala 77:18:@284.6]
  assign _GEN_103 = 3'h5 == _T_1158 ? 1'h0 : _GEN_102; // @[StoreQueue.scala 77:18:@284.6]
  assign _GEN_104 = 3'h6 == _T_1158 ? 1'h0 : _GEN_103; // @[StoreQueue.scala 77:18:@284.6]
  assign _GEN_105 = 3'h7 == _T_1158 ? 1'h0 : _GEN_104; // @[StoreQueue.scala 77:18:@284.6]
  assign _GEN_106 = initBits_5 ? _GEN_97 : offsetQ_5; // @[StoreQueue.scala 75:25:@270.4]
  assign _GEN_107 = initBits_5 ? _GEN_105 : portQ_5; // @[StoreQueue.scala 75:25:@270.4]
  assign _T_1176 = _T_1013[2:0]; // @[:@292.6]
  assign _GEN_109 = 3'h1 == _T_1176 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_110 = 3'h2 == _T_1176 ? io_bbStoreOffsets_2 : _GEN_109; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_111 = 3'h3 == _T_1176 ? io_bbStoreOffsets_3 : _GEN_110; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_112 = 3'h4 == _T_1176 ? io_bbStoreOffsets_4 : _GEN_111; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_113 = 3'h5 == _T_1176 ? io_bbStoreOffsets_5 : _GEN_112; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_114 = 3'h6 == _T_1176 ? io_bbStoreOffsets_6 : _GEN_113; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_115 = 3'h7 == _T_1176 ? io_bbStoreOffsets_7 : _GEN_114; // @[StoreQueue.scala 76:20:@293.6]
  assign _GEN_117 = 3'h1 == _T_1176 ? io_bbStorePorts_1 : 1'h0; // @[StoreQueue.scala 77:18:@300.6]
  assign _GEN_118 = 3'h2 == _T_1176 ? 1'h0 : _GEN_117; // @[StoreQueue.scala 77:18:@300.6]
  assign _GEN_119 = 3'h3 == _T_1176 ? 1'h0 : _GEN_118; // @[StoreQueue.scala 77:18:@300.6]
  assign _GEN_120 = 3'h4 == _T_1176 ? 1'h0 : _GEN_119; // @[StoreQueue.scala 77:18:@300.6]
  assign _GEN_121 = 3'h5 == _T_1176 ? 1'h0 : _GEN_120; // @[StoreQueue.scala 77:18:@300.6]
  assign _GEN_122 = 3'h6 == _T_1176 ? 1'h0 : _GEN_121; // @[StoreQueue.scala 77:18:@300.6]
  assign _GEN_123 = 3'h7 == _T_1176 ? 1'h0 : _GEN_122; // @[StoreQueue.scala 77:18:@300.6]
  assign _GEN_124 = initBits_6 ? _GEN_115 : offsetQ_6; // @[StoreQueue.scala 75:25:@286.4]
  assign _GEN_125 = initBits_6 ? _GEN_123 : portQ_6; // @[StoreQueue.scala 75:25:@286.4]
  assign _T_1194 = _T_1022[2:0]; // @[:@308.6]
  assign _GEN_127 = 3'h1 == _T_1194 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_128 = 3'h2 == _T_1194 ? io_bbStoreOffsets_2 : _GEN_127; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_129 = 3'h3 == _T_1194 ? io_bbStoreOffsets_3 : _GEN_128; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_130 = 3'h4 == _T_1194 ? io_bbStoreOffsets_4 : _GEN_129; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_131 = 3'h5 == _T_1194 ? io_bbStoreOffsets_5 : _GEN_130; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_132 = 3'h6 == _T_1194 ? io_bbStoreOffsets_6 : _GEN_131; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_133 = 3'h7 == _T_1194 ? io_bbStoreOffsets_7 : _GEN_132; // @[StoreQueue.scala 76:20:@309.6]
  assign _GEN_135 = 3'h1 == _T_1194 ? io_bbStorePorts_1 : 1'h0; // @[StoreQueue.scala 77:18:@316.6]
  assign _GEN_136 = 3'h2 == _T_1194 ? 1'h0 : _GEN_135; // @[StoreQueue.scala 77:18:@316.6]
  assign _GEN_137 = 3'h3 == _T_1194 ? 1'h0 : _GEN_136; // @[StoreQueue.scala 77:18:@316.6]
  assign _GEN_138 = 3'h4 == _T_1194 ? 1'h0 : _GEN_137; // @[StoreQueue.scala 77:18:@316.6]
  assign _GEN_139 = 3'h5 == _T_1194 ? 1'h0 : _GEN_138; // @[StoreQueue.scala 77:18:@316.6]
  assign _GEN_140 = 3'h6 == _T_1194 ? 1'h0 : _GEN_139; // @[StoreQueue.scala 77:18:@316.6]
  assign _GEN_141 = 3'h7 == _T_1194 ? 1'h0 : _GEN_140; // @[StoreQueue.scala 77:18:@316.6]
  assign _GEN_142 = initBits_7 ? _GEN_133 : offsetQ_7; // @[StoreQueue.scala 75:25:@302.4]
  assign _GEN_143 = initBits_7 ? _GEN_141 : portQ_7; // @[StoreQueue.scala 75:25:@302.4]
  assign _T_1216 = _GEN_7 + 3'h1; // @[util.scala 10:8:@327.6]
  assign _GEN_72 = _T_1216 % 4'h8; // @[util.scala 10:14:@328.6]
  assign _T_1217 = _GEN_72[3:0]; // @[util.scala 10:14:@328.6]
  assign _GEN_443 = {{1'd0}, io_loadTail}; // @[StoreQueue.scala 96:56:@329.6]
  assign _T_1218 = _T_1217 == _GEN_443; // @[StoreQueue.scala 96:56:@329.6]
  assign _T_1219 = io_loadEmpty & _T_1218; // @[StoreQueue.scala 95:50:@330.6]
  assign _T_1221 = _T_1219 == 1'h0; // @[StoreQueue.scala 95:35:@331.6]
  assign _T_1223 = previousLoadHead <= offsetQ_0; // @[StoreQueue.scala 100:35:@339.8]
  assign _T_1224 = offsetQ_0 < io_loadHead; // @[StoreQueue.scala 100:87:@340.8]
  assign _T_1225 = _T_1223 & _T_1224; // @[StoreQueue.scala 100:61:@341.8]
  assign _T_1227 = previousLoadHead > io_loadHead; // @[StoreQueue.scala 102:35:@346.10]
  assign _T_1228 = io_loadHead <= offsetQ_0; // @[StoreQueue.scala 103:23:@347.10]
  assign _T_1229 = offsetQ_0 < previousLoadHead; // @[StoreQueue.scala 103:75:@348.10]
  assign _T_1230 = _T_1228 & _T_1229; // @[StoreQueue.scala 103:49:@349.10]
  assign _T_1232 = _T_1230 == 1'h0; // @[StoreQueue.scala 103:9:@350.10]
  assign _T_1233 = _T_1227 & _T_1232; // @[StoreQueue.scala 102:49:@351.10]
  assign _GEN_152 = _T_1233 ? 1'h0 : checkBits_0; // @[StoreQueue.scala 103:96:@352.10]
  assign _GEN_153 = _T_1225 ? 1'h0 : _GEN_152; // @[StoreQueue.scala 100:102:@342.8]
  assign _GEN_154 = io_loadEmpty ? 1'h0 : _GEN_153; // @[StoreQueue.scala 98:26:@335.6]
  assign _GEN_155 = initBits_0 ? _T_1221 : _GEN_154; // @[StoreQueue.scala 94:35:@320.4]
  assign _T_1246 = _GEN_25 + 3'h1; // @[util.scala 10:8:@363.6]
  assign _GEN_80 = _T_1246 % 4'h8; // @[util.scala 10:14:@364.6]
  assign _T_1247 = _GEN_80[3:0]; // @[util.scala 10:14:@364.6]
  assign _T_1248 = _T_1247 == _GEN_443; // @[StoreQueue.scala 96:56:@365.6]
  assign _T_1249 = io_loadEmpty & _T_1248; // @[StoreQueue.scala 95:50:@366.6]
  assign _T_1251 = _T_1249 == 1'h0; // @[StoreQueue.scala 95:35:@367.6]
  assign _T_1253 = previousLoadHead <= offsetQ_1; // @[StoreQueue.scala 100:35:@375.8]
  assign _T_1254 = offsetQ_1 < io_loadHead; // @[StoreQueue.scala 100:87:@376.8]
  assign _T_1255 = _T_1253 & _T_1254; // @[StoreQueue.scala 100:61:@377.8]
  assign _T_1258 = io_loadHead <= offsetQ_1; // @[StoreQueue.scala 103:23:@383.10]
  assign _T_1259 = offsetQ_1 < previousLoadHead; // @[StoreQueue.scala 103:75:@384.10]
  assign _T_1260 = _T_1258 & _T_1259; // @[StoreQueue.scala 103:49:@385.10]
  assign _T_1262 = _T_1260 == 1'h0; // @[StoreQueue.scala 103:9:@386.10]
  assign _T_1263 = _T_1227 & _T_1262; // @[StoreQueue.scala 102:49:@387.10]
  assign _GEN_164 = _T_1263 ? 1'h0 : checkBits_1; // @[StoreQueue.scala 103:96:@388.10]
  assign _GEN_165 = _T_1255 ? 1'h0 : _GEN_164; // @[StoreQueue.scala 100:102:@378.8]
  assign _GEN_166 = io_loadEmpty ? 1'h0 : _GEN_165; // @[StoreQueue.scala 98:26:@371.6]
  assign _GEN_167 = initBits_1 ? _T_1251 : _GEN_166; // @[StoreQueue.scala 94:35:@356.4]
  assign _T_1276 = _GEN_43 + 3'h1; // @[util.scala 10:8:@399.6]
  assign _GEN_90 = _T_1276 % 4'h8; // @[util.scala 10:14:@400.6]
  assign _T_1277 = _GEN_90[3:0]; // @[util.scala 10:14:@400.6]
  assign _T_1278 = _T_1277 == _GEN_443; // @[StoreQueue.scala 96:56:@401.6]
  assign _T_1279 = io_loadEmpty & _T_1278; // @[StoreQueue.scala 95:50:@402.6]
  assign _T_1281 = _T_1279 == 1'h0; // @[StoreQueue.scala 95:35:@403.6]
  assign _T_1283 = previousLoadHead <= offsetQ_2; // @[StoreQueue.scala 100:35:@411.8]
  assign _T_1284 = offsetQ_2 < io_loadHead; // @[StoreQueue.scala 100:87:@412.8]
  assign _T_1285 = _T_1283 & _T_1284; // @[StoreQueue.scala 100:61:@413.8]
  assign _T_1288 = io_loadHead <= offsetQ_2; // @[StoreQueue.scala 103:23:@419.10]
  assign _T_1289 = offsetQ_2 < previousLoadHead; // @[StoreQueue.scala 103:75:@420.10]
  assign _T_1290 = _T_1288 & _T_1289; // @[StoreQueue.scala 103:49:@421.10]
  assign _T_1292 = _T_1290 == 1'h0; // @[StoreQueue.scala 103:9:@422.10]
  assign _T_1293 = _T_1227 & _T_1292; // @[StoreQueue.scala 102:49:@423.10]
  assign _GEN_176 = _T_1293 ? 1'h0 : checkBits_2; // @[StoreQueue.scala 103:96:@424.10]
  assign _GEN_177 = _T_1285 ? 1'h0 : _GEN_176; // @[StoreQueue.scala 100:102:@414.8]
  assign _GEN_178 = io_loadEmpty ? 1'h0 : _GEN_177; // @[StoreQueue.scala 98:26:@407.6]
  assign _GEN_179 = initBits_2 ? _T_1281 : _GEN_178; // @[StoreQueue.scala 94:35:@392.4]
  assign _T_1306 = _GEN_61 + 3'h1; // @[util.scala 10:8:@435.6]
  assign _GEN_98 = _T_1306 % 4'h8; // @[util.scala 10:14:@436.6]
  assign _T_1307 = _GEN_98[3:0]; // @[util.scala 10:14:@436.6]
  assign _T_1308 = _T_1307 == _GEN_443; // @[StoreQueue.scala 96:56:@437.6]
  assign _T_1309 = io_loadEmpty & _T_1308; // @[StoreQueue.scala 95:50:@438.6]
  assign _T_1311 = _T_1309 == 1'h0; // @[StoreQueue.scala 95:35:@439.6]
  assign _T_1313 = previousLoadHead <= offsetQ_3; // @[StoreQueue.scala 100:35:@447.8]
  assign _T_1314 = offsetQ_3 < io_loadHead; // @[StoreQueue.scala 100:87:@448.8]
  assign _T_1315 = _T_1313 & _T_1314; // @[StoreQueue.scala 100:61:@449.8]
  assign _T_1318 = io_loadHead <= offsetQ_3; // @[StoreQueue.scala 103:23:@455.10]
  assign _T_1319 = offsetQ_3 < previousLoadHead; // @[StoreQueue.scala 103:75:@456.10]
  assign _T_1320 = _T_1318 & _T_1319; // @[StoreQueue.scala 103:49:@457.10]
  assign _T_1322 = _T_1320 == 1'h0; // @[StoreQueue.scala 103:9:@458.10]
  assign _T_1323 = _T_1227 & _T_1322; // @[StoreQueue.scala 102:49:@459.10]
  assign _GEN_188 = _T_1323 ? 1'h0 : checkBits_3; // @[StoreQueue.scala 103:96:@460.10]
  assign _GEN_189 = _T_1315 ? 1'h0 : _GEN_188; // @[StoreQueue.scala 100:102:@450.8]
  assign _GEN_190 = io_loadEmpty ? 1'h0 : _GEN_189; // @[StoreQueue.scala 98:26:@443.6]
  assign _GEN_191 = initBits_3 ? _T_1311 : _GEN_190; // @[StoreQueue.scala 94:35:@428.4]
  assign _T_1336 = _GEN_79 + 3'h1; // @[util.scala 10:8:@471.6]
  assign _GEN_108 = _T_1336 % 4'h8; // @[util.scala 10:14:@472.6]
  assign _T_1337 = _GEN_108[3:0]; // @[util.scala 10:14:@472.6]
  assign _T_1338 = _T_1337 == _GEN_443; // @[StoreQueue.scala 96:56:@473.6]
  assign _T_1339 = io_loadEmpty & _T_1338; // @[StoreQueue.scala 95:50:@474.6]
  assign _T_1341 = _T_1339 == 1'h0; // @[StoreQueue.scala 95:35:@475.6]
  assign _T_1343 = previousLoadHead <= offsetQ_4; // @[StoreQueue.scala 100:35:@483.8]
  assign _T_1344 = offsetQ_4 < io_loadHead; // @[StoreQueue.scala 100:87:@484.8]
  assign _T_1345 = _T_1343 & _T_1344; // @[StoreQueue.scala 100:61:@485.8]
  assign _T_1348 = io_loadHead <= offsetQ_4; // @[StoreQueue.scala 103:23:@491.10]
  assign _T_1349 = offsetQ_4 < previousLoadHead; // @[StoreQueue.scala 103:75:@492.10]
  assign _T_1350 = _T_1348 & _T_1349; // @[StoreQueue.scala 103:49:@493.10]
  assign _T_1352 = _T_1350 == 1'h0; // @[StoreQueue.scala 103:9:@494.10]
  assign _T_1353 = _T_1227 & _T_1352; // @[StoreQueue.scala 102:49:@495.10]
  assign _GEN_200 = _T_1353 ? 1'h0 : checkBits_4; // @[StoreQueue.scala 103:96:@496.10]
  assign _GEN_201 = _T_1345 ? 1'h0 : _GEN_200; // @[StoreQueue.scala 100:102:@486.8]
  assign _GEN_202 = io_loadEmpty ? 1'h0 : _GEN_201; // @[StoreQueue.scala 98:26:@479.6]
  assign _GEN_203 = initBits_4 ? _T_1341 : _GEN_202; // @[StoreQueue.scala 94:35:@464.4]
  assign _T_1366 = _GEN_97 + 3'h1; // @[util.scala 10:8:@507.6]
  assign _GEN_116 = _T_1366 % 4'h8; // @[util.scala 10:14:@508.6]
  assign _T_1367 = _GEN_116[3:0]; // @[util.scala 10:14:@508.6]
  assign _T_1368 = _T_1367 == _GEN_443; // @[StoreQueue.scala 96:56:@509.6]
  assign _T_1369 = io_loadEmpty & _T_1368; // @[StoreQueue.scala 95:50:@510.6]
  assign _T_1371 = _T_1369 == 1'h0; // @[StoreQueue.scala 95:35:@511.6]
  assign _T_1373 = previousLoadHead <= offsetQ_5; // @[StoreQueue.scala 100:35:@519.8]
  assign _T_1374 = offsetQ_5 < io_loadHead; // @[StoreQueue.scala 100:87:@520.8]
  assign _T_1375 = _T_1373 & _T_1374; // @[StoreQueue.scala 100:61:@521.8]
  assign _T_1378 = io_loadHead <= offsetQ_5; // @[StoreQueue.scala 103:23:@527.10]
  assign _T_1379 = offsetQ_5 < previousLoadHead; // @[StoreQueue.scala 103:75:@528.10]
  assign _T_1380 = _T_1378 & _T_1379; // @[StoreQueue.scala 103:49:@529.10]
  assign _T_1382 = _T_1380 == 1'h0; // @[StoreQueue.scala 103:9:@530.10]
  assign _T_1383 = _T_1227 & _T_1382; // @[StoreQueue.scala 102:49:@531.10]
  assign _GEN_212 = _T_1383 ? 1'h0 : checkBits_5; // @[StoreQueue.scala 103:96:@532.10]
  assign _GEN_213 = _T_1375 ? 1'h0 : _GEN_212; // @[StoreQueue.scala 100:102:@522.8]
  assign _GEN_214 = io_loadEmpty ? 1'h0 : _GEN_213; // @[StoreQueue.scala 98:26:@515.6]
  assign _GEN_215 = initBits_5 ? _T_1371 : _GEN_214; // @[StoreQueue.scala 94:35:@500.4]
  assign _T_1396 = _GEN_115 + 3'h1; // @[util.scala 10:8:@543.6]
  assign _GEN_126 = _T_1396 % 4'h8; // @[util.scala 10:14:@544.6]
  assign _T_1397 = _GEN_126[3:0]; // @[util.scala 10:14:@544.6]
  assign _T_1398 = _T_1397 == _GEN_443; // @[StoreQueue.scala 96:56:@545.6]
  assign _T_1399 = io_loadEmpty & _T_1398; // @[StoreQueue.scala 95:50:@546.6]
  assign _T_1401 = _T_1399 == 1'h0; // @[StoreQueue.scala 95:35:@547.6]
  assign _T_1403 = previousLoadHead <= offsetQ_6; // @[StoreQueue.scala 100:35:@555.8]
  assign _T_1404 = offsetQ_6 < io_loadHead; // @[StoreQueue.scala 100:87:@556.8]
  assign _T_1405 = _T_1403 & _T_1404; // @[StoreQueue.scala 100:61:@557.8]
  assign _T_1408 = io_loadHead <= offsetQ_6; // @[StoreQueue.scala 103:23:@563.10]
  assign _T_1409 = offsetQ_6 < previousLoadHead; // @[StoreQueue.scala 103:75:@564.10]
  assign _T_1410 = _T_1408 & _T_1409; // @[StoreQueue.scala 103:49:@565.10]
  assign _T_1412 = _T_1410 == 1'h0; // @[StoreQueue.scala 103:9:@566.10]
  assign _T_1413 = _T_1227 & _T_1412; // @[StoreQueue.scala 102:49:@567.10]
  assign _GEN_224 = _T_1413 ? 1'h0 : checkBits_6; // @[StoreQueue.scala 103:96:@568.10]
  assign _GEN_225 = _T_1405 ? 1'h0 : _GEN_224; // @[StoreQueue.scala 100:102:@558.8]
  assign _GEN_226 = io_loadEmpty ? 1'h0 : _GEN_225; // @[StoreQueue.scala 98:26:@551.6]
  assign _GEN_227 = initBits_6 ? _T_1401 : _GEN_226; // @[StoreQueue.scala 94:35:@536.4]
  assign _T_1426 = _GEN_133 + 3'h1; // @[util.scala 10:8:@579.6]
  assign _GEN_134 = _T_1426 % 4'h8; // @[util.scala 10:14:@580.6]
  assign _T_1427 = _GEN_134[3:0]; // @[util.scala 10:14:@580.6]
  assign _T_1428 = _T_1427 == _GEN_443; // @[StoreQueue.scala 96:56:@581.6]
  assign _T_1429 = io_loadEmpty & _T_1428; // @[StoreQueue.scala 95:50:@582.6]
  assign _T_1431 = _T_1429 == 1'h0; // @[StoreQueue.scala 95:35:@583.6]
  assign _T_1433 = previousLoadHead <= offsetQ_7; // @[StoreQueue.scala 100:35:@591.8]
  assign _T_1434 = offsetQ_7 < io_loadHead; // @[StoreQueue.scala 100:87:@592.8]
  assign _T_1435 = _T_1433 & _T_1434; // @[StoreQueue.scala 100:61:@593.8]
  assign _T_1438 = io_loadHead <= offsetQ_7; // @[StoreQueue.scala 103:23:@599.10]
  assign _T_1439 = offsetQ_7 < previousLoadHead; // @[StoreQueue.scala 103:75:@600.10]
  assign _T_1440 = _T_1438 & _T_1439; // @[StoreQueue.scala 103:49:@601.10]
  assign _T_1442 = _T_1440 == 1'h0; // @[StoreQueue.scala 103:9:@602.10]
  assign _T_1443 = _T_1227 & _T_1442; // @[StoreQueue.scala 102:49:@603.10]
  assign _GEN_236 = _T_1443 ? 1'h0 : checkBits_7; // @[StoreQueue.scala 103:96:@604.10]
  assign _GEN_237 = _T_1435 ? 1'h0 : _GEN_236; // @[StoreQueue.scala 100:102:@594.8]
  assign _GEN_238 = io_loadEmpty ? 1'h0 : _GEN_237; // @[StoreQueue.scala 98:26:@587.6]
  assign _GEN_239 = initBits_7 ? _T_1431 : _GEN_238; // @[StoreQueue.scala 94:35:@572.4]
  assign _T_1445 = io_loadHead < io_loadTail; // @[StoreQueue.scala 119:103:@608.4]
  assign _T_1447 = io_loadHead <= 3'h0; // @[StoreQueue.scala 120:17:@609.4]
  assign _T_1449 = 3'h0 < io_loadTail; // @[StoreQueue.scala 120:35:@610.4]
  assign _T_1450 = _T_1447 & _T_1449; // @[StoreQueue.scala 120:26:@611.4]
  assign _T_1452 = io_loadEmpty == 1'h0; // @[StoreQueue.scala 120:50:@612.4]
  assign _T_1454 = io_loadTail <= 3'h0; // @[StoreQueue.scala 120:81:@613.4]
  assign _T_1456 = 3'h0 < io_loadHead; // @[StoreQueue.scala 120:99:@614.4]
  assign _T_1457 = _T_1454 & _T_1456; // @[StoreQueue.scala 120:90:@615.4]
  assign _T_1459 = _T_1457 == 1'h0; // @[StoreQueue.scala 120:67:@616.4]
  assign _T_1460 = _T_1452 & _T_1459; // @[StoreQueue.scala 120:64:@617.4]
  assign validEntriesInLoadQ_0 = _T_1445 ? _T_1450 : _T_1460; // @[StoreQueue.scala 119:90:@618.4]
  assign _T_1464 = io_loadHead <= 3'h1; // @[StoreQueue.scala 120:17:@620.4]
  assign _T_1466 = 3'h1 < io_loadTail; // @[StoreQueue.scala 120:35:@621.4]
  assign _T_1467 = _T_1464 & _T_1466; // @[StoreQueue.scala 120:26:@622.4]
  assign _T_1471 = io_loadTail <= 3'h1; // @[StoreQueue.scala 120:81:@624.4]
  assign _T_1473 = 3'h1 < io_loadHead; // @[StoreQueue.scala 120:99:@625.4]
  assign _T_1474 = _T_1471 & _T_1473; // @[StoreQueue.scala 120:90:@626.4]
  assign _T_1476 = _T_1474 == 1'h0; // @[StoreQueue.scala 120:67:@627.4]
  assign _T_1477 = _T_1452 & _T_1476; // @[StoreQueue.scala 120:64:@628.4]
  assign validEntriesInLoadQ_1 = _T_1445 ? _T_1467 : _T_1477; // @[StoreQueue.scala 119:90:@629.4]
  assign _T_1481 = io_loadHead <= 3'h2; // @[StoreQueue.scala 120:17:@631.4]
  assign _T_1483 = 3'h2 < io_loadTail; // @[StoreQueue.scala 120:35:@632.4]
  assign _T_1484 = _T_1481 & _T_1483; // @[StoreQueue.scala 120:26:@633.4]
  assign _T_1488 = io_loadTail <= 3'h2; // @[StoreQueue.scala 120:81:@635.4]
  assign _T_1490 = 3'h2 < io_loadHead; // @[StoreQueue.scala 120:99:@636.4]
  assign _T_1491 = _T_1488 & _T_1490; // @[StoreQueue.scala 120:90:@637.4]
  assign _T_1493 = _T_1491 == 1'h0; // @[StoreQueue.scala 120:67:@638.4]
  assign _T_1494 = _T_1452 & _T_1493; // @[StoreQueue.scala 120:64:@639.4]
  assign validEntriesInLoadQ_2 = _T_1445 ? _T_1484 : _T_1494; // @[StoreQueue.scala 119:90:@640.4]
  assign _T_1498 = io_loadHead <= 3'h3; // @[StoreQueue.scala 120:17:@642.4]
  assign _T_1500 = 3'h3 < io_loadTail; // @[StoreQueue.scala 120:35:@643.4]
  assign _T_1501 = _T_1498 & _T_1500; // @[StoreQueue.scala 120:26:@644.4]
  assign _T_1505 = io_loadTail <= 3'h3; // @[StoreQueue.scala 120:81:@646.4]
  assign _T_1507 = 3'h3 < io_loadHead; // @[StoreQueue.scala 120:99:@647.4]
  assign _T_1508 = _T_1505 & _T_1507; // @[StoreQueue.scala 120:90:@648.4]
  assign _T_1510 = _T_1508 == 1'h0; // @[StoreQueue.scala 120:67:@649.4]
  assign _T_1511 = _T_1452 & _T_1510; // @[StoreQueue.scala 120:64:@650.4]
  assign validEntriesInLoadQ_3 = _T_1445 ? _T_1501 : _T_1511; // @[StoreQueue.scala 119:90:@651.4]
  assign _T_1515 = io_loadHead <= 3'h4; // @[StoreQueue.scala 120:17:@653.4]
  assign _T_1517 = 3'h4 < io_loadTail; // @[StoreQueue.scala 120:35:@654.4]
  assign _T_1518 = _T_1515 & _T_1517; // @[StoreQueue.scala 120:26:@655.4]
  assign _T_1522 = io_loadTail <= 3'h4; // @[StoreQueue.scala 120:81:@657.4]
  assign _T_1524 = 3'h4 < io_loadHead; // @[StoreQueue.scala 120:99:@658.4]
  assign _T_1525 = _T_1522 & _T_1524; // @[StoreQueue.scala 120:90:@659.4]
  assign _T_1527 = _T_1525 == 1'h0; // @[StoreQueue.scala 120:67:@660.4]
  assign _T_1528 = _T_1452 & _T_1527; // @[StoreQueue.scala 120:64:@661.4]
  assign validEntriesInLoadQ_4 = _T_1445 ? _T_1518 : _T_1528; // @[StoreQueue.scala 119:90:@662.4]
  assign _T_1532 = io_loadHead <= 3'h5; // @[StoreQueue.scala 120:17:@664.4]
  assign _T_1534 = 3'h5 < io_loadTail; // @[StoreQueue.scala 120:35:@665.4]
  assign _T_1535 = _T_1532 & _T_1534; // @[StoreQueue.scala 120:26:@666.4]
  assign _T_1539 = io_loadTail <= 3'h5; // @[StoreQueue.scala 120:81:@668.4]
  assign _T_1541 = 3'h5 < io_loadHead; // @[StoreQueue.scala 120:99:@669.4]
  assign _T_1542 = _T_1539 & _T_1541; // @[StoreQueue.scala 120:90:@670.4]
  assign _T_1544 = _T_1542 == 1'h0; // @[StoreQueue.scala 120:67:@671.4]
  assign _T_1545 = _T_1452 & _T_1544; // @[StoreQueue.scala 120:64:@672.4]
  assign validEntriesInLoadQ_5 = _T_1445 ? _T_1535 : _T_1545; // @[StoreQueue.scala 119:90:@673.4]
  assign _T_1549 = io_loadHead <= 3'h6; // @[StoreQueue.scala 120:17:@675.4]
  assign _T_1551 = 3'h6 < io_loadTail; // @[StoreQueue.scala 120:35:@676.4]
  assign _T_1552 = _T_1549 & _T_1551; // @[StoreQueue.scala 120:26:@677.4]
  assign _T_1556 = io_loadTail <= 3'h6; // @[StoreQueue.scala 120:81:@679.4]
  assign _T_1558 = 3'h6 < io_loadHead; // @[StoreQueue.scala 120:99:@680.4]
  assign _T_1559 = _T_1556 & _T_1558; // @[StoreQueue.scala 120:90:@681.4]
  assign _T_1561 = _T_1559 == 1'h0; // @[StoreQueue.scala 120:67:@682.4]
  assign _T_1562 = _T_1452 & _T_1561; // @[StoreQueue.scala 120:64:@683.4]
  assign validEntriesInLoadQ_6 = _T_1445 ? _T_1552 : _T_1562; // @[StoreQueue.scala 119:90:@684.4]
  assign validEntriesInLoadQ_7 = _T_1445 ? 1'h0 : _T_1452; // @[StoreQueue.scala 119:90:@695.4]
  assign _GEN_241 = 3'h1 == head ? offsetQ_1 : offsetQ_0; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_242 = 3'h2 == head ? offsetQ_2 : _GEN_241; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_243 = 3'h3 == head ? offsetQ_3 : _GEN_242; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_244 = 3'h4 == head ? offsetQ_4 : _GEN_243; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_245 = 3'h5 == head ? offsetQ_5 : _GEN_244; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_246 = 3'h6 == head ? offsetQ_6 : _GEN_245; // @[StoreQueue.scala 126:96:@705.4]
  assign _GEN_247 = 3'h7 == head ? offsetQ_7 : _GEN_246; // @[StoreQueue.scala 126:96:@705.4]
  assign _T_1597 = io_loadHead <= _GEN_247; // @[StoreQueue.scala 126:96:@705.4]
  assign loadsToCheck_0 = _T_1597 ? _T_1447 : 1'h1; // @[StoreQueue.scala 126:83:@713.4]
  assign _T_1627 = 3'h1 <= _GEN_247; // @[StoreQueue.scala 127:37:@716.4]
  assign _T_1628 = _T_1464 & _T_1627; // @[StoreQueue.scala 127:28:@717.4]
  assign _T_1633 = _GEN_247 < 3'h1; // @[StoreQueue.scala 127:71:@718.4]
  assign _T_1636 = _T_1633 & _T_1473; // @[StoreQueue.scala 127:79:@720.4]
  assign _T_1638 = _T_1636 == 1'h0; // @[StoreQueue.scala 127:55:@721.4]
  assign loadsToCheck_1 = _T_1597 ? _T_1628 : _T_1638; // @[StoreQueue.scala 126:83:@722.4]
  assign _T_1650 = 3'h2 <= _GEN_247; // @[StoreQueue.scala 127:37:@725.4]
  assign _T_1651 = _T_1481 & _T_1650; // @[StoreQueue.scala 127:28:@726.4]
  assign _T_1656 = _GEN_247 < 3'h2; // @[StoreQueue.scala 127:71:@727.4]
  assign _T_1659 = _T_1656 & _T_1490; // @[StoreQueue.scala 127:79:@729.4]
  assign _T_1661 = _T_1659 == 1'h0; // @[StoreQueue.scala 127:55:@730.4]
  assign loadsToCheck_2 = _T_1597 ? _T_1651 : _T_1661; // @[StoreQueue.scala 126:83:@731.4]
  assign _T_1673 = 3'h3 <= _GEN_247; // @[StoreQueue.scala 127:37:@734.4]
  assign _T_1674 = _T_1498 & _T_1673; // @[StoreQueue.scala 127:28:@735.4]
  assign _T_1679 = _GEN_247 < 3'h3; // @[StoreQueue.scala 127:71:@736.4]
  assign _T_1682 = _T_1679 & _T_1507; // @[StoreQueue.scala 127:79:@738.4]
  assign _T_1684 = _T_1682 == 1'h0; // @[StoreQueue.scala 127:55:@739.4]
  assign loadsToCheck_3 = _T_1597 ? _T_1674 : _T_1684; // @[StoreQueue.scala 126:83:@740.4]
  assign _T_1696 = 3'h4 <= _GEN_247; // @[StoreQueue.scala 127:37:@743.4]
  assign _T_1697 = _T_1515 & _T_1696; // @[StoreQueue.scala 127:28:@744.4]
  assign _T_1702 = _GEN_247 < 3'h4; // @[StoreQueue.scala 127:71:@745.4]
  assign _T_1705 = _T_1702 & _T_1524; // @[StoreQueue.scala 127:79:@747.4]
  assign _T_1707 = _T_1705 == 1'h0; // @[StoreQueue.scala 127:55:@748.4]
  assign loadsToCheck_4 = _T_1597 ? _T_1697 : _T_1707; // @[StoreQueue.scala 126:83:@749.4]
  assign _T_1719 = 3'h5 <= _GEN_247; // @[StoreQueue.scala 127:37:@752.4]
  assign _T_1720 = _T_1532 & _T_1719; // @[StoreQueue.scala 127:28:@753.4]
  assign _T_1725 = _GEN_247 < 3'h5; // @[StoreQueue.scala 127:71:@754.4]
  assign _T_1728 = _T_1725 & _T_1541; // @[StoreQueue.scala 127:79:@756.4]
  assign _T_1730 = _T_1728 == 1'h0; // @[StoreQueue.scala 127:55:@757.4]
  assign loadsToCheck_5 = _T_1597 ? _T_1720 : _T_1730; // @[StoreQueue.scala 126:83:@758.4]
  assign _T_1742 = 3'h6 <= _GEN_247; // @[StoreQueue.scala 127:37:@761.4]
  assign _T_1743 = _T_1549 & _T_1742; // @[StoreQueue.scala 127:28:@762.4]
  assign _T_1748 = _GEN_247 < 3'h6; // @[StoreQueue.scala 127:71:@763.4]
  assign _T_1751 = _T_1748 & _T_1558; // @[StoreQueue.scala 127:79:@765.4]
  assign _T_1753 = _T_1751 == 1'h0; // @[StoreQueue.scala 127:55:@766.4]
  assign loadsToCheck_6 = _T_1597 ? _T_1743 : _T_1753; // @[StoreQueue.scala 126:83:@767.4]
  assign _T_1765 = 3'h7 <= _GEN_247; // @[StoreQueue.scala 127:37:@770.4]
  assign loadsToCheck_7 = _T_1597 ? _T_1765 : 1'h1; // @[StoreQueue.scala 126:83:@776.4]
  assign _T_1791 = loadsToCheck_0 & validEntriesInLoadQ_0; // @[StoreQueue.scala 133:16:@786.4]
  assign _GEN_249 = 3'h1 == head ? checkBits_1 : checkBits_0; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_250 = 3'h2 == head ? checkBits_2 : _GEN_249; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_251 = 3'h3 == head ? checkBits_3 : _GEN_250; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_252 = 3'h4 == head ? checkBits_4 : _GEN_251; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_253 = 3'h5 == head ? checkBits_5 : _GEN_252; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_254 = 3'h6 == head ? checkBits_6 : _GEN_253; // @[StoreQueue.scala 133:24:@787.4]
  assign _GEN_255 = 3'h7 == head ? checkBits_7 : _GEN_254; // @[StoreQueue.scala 133:24:@787.4]
  assign entriesToCheck_0 = _T_1791 & _GEN_255; // @[StoreQueue.scala 133:24:@787.4]
  assign _T_1796 = loadsToCheck_1 & validEntriesInLoadQ_1; // @[StoreQueue.scala 133:16:@788.4]
  assign entriesToCheck_1 = _T_1796 & _GEN_255; // @[StoreQueue.scala 133:24:@789.4]
  assign _T_1801 = loadsToCheck_2 & validEntriesInLoadQ_2; // @[StoreQueue.scala 133:16:@790.4]
  assign entriesToCheck_2 = _T_1801 & _GEN_255; // @[StoreQueue.scala 133:24:@791.4]
  assign _T_1806 = loadsToCheck_3 & validEntriesInLoadQ_3; // @[StoreQueue.scala 133:16:@792.4]
  assign entriesToCheck_3 = _T_1806 & _GEN_255; // @[StoreQueue.scala 133:24:@793.4]
  assign _T_1811 = loadsToCheck_4 & validEntriesInLoadQ_4; // @[StoreQueue.scala 133:16:@794.4]
  assign entriesToCheck_4 = _T_1811 & _GEN_255; // @[StoreQueue.scala 133:24:@795.4]
  assign _T_1816 = loadsToCheck_5 & validEntriesInLoadQ_5; // @[StoreQueue.scala 133:16:@796.4]
  assign entriesToCheck_5 = _T_1816 & _GEN_255; // @[StoreQueue.scala 133:24:@797.4]
  assign _T_1821 = loadsToCheck_6 & validEntriesInLoadQ_6; // @[StoreQueue.scala 133:16:@798.4]
  assign entriesToCheck_6 = _T_1821 & _GEN_255; // @[StoreQueue.scala 133:24:@799.4]
  assign _T_1826 = loadsToCheck_7 & validEntriesInLoadQ_7; // @[StoreQueue.scala 133:16:@800.4]
  assign entriesToCheck_7 = _T_1826 & _GEN_255; // @[StoreQueue.scala 133:24:@801.4]
  assign _T_1858 = entriesToCheck_0 == 1'h0; // @[StoreQueue.scala 140:34:@812.4]
  assign _T_1859 = _T_1858 | io_loadDataDone_0; // @[StoreQueue.scala 140:64:@813.4]
  assign _GEN_257 = 3'h1 == head ? addrQ_1 : addrQ_0; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_258 = 3'h2 == head ? addrQ_2 : _GEN_257; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_259 = 3'h3 == head ? addrQ_3 : _GEN_258; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_260 = 3'h4 == head ? addrQ_4 : _GEN_259; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_261 = 3'h5 == head ? addrQ_5 : _GEN_260; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_262 = 3'h6 == head ? addrQ_6 : _GEN_261; // @[StoreQueue.scala 141:51:@814.4]
  assign _GEN_263 = 3'h7 == head ? addrQ_7 : _GEN_262; // @[StoreQueue.scala 141:51:@814.4]
  assign _T_1863 = _GEN_263 != io_loadAddressQueue_0; // @[StoreQueue.scala 141:51:@814.4]
  assign _T_1864 = io_loadAddressDone_0 & _T_1863; // @[StoreQueue.scala 141:36:@815.4]
  assign noConflicts_0 = _T_1859 | _T_1864; // @[StoreQueue.scala 140:95:@816.4]
  assign _T_1867 = entriesToCheck_1 == 1'h0; // @[StoreQueue.scala 140:34:@818.4]
  assign _T_1868 = _T_1867 | io_loadDataDone_1; // @[StoreQueue.scala 140:64:@819.4]
  assign _T_1872 = _GEN_263 != io_loadAddressQueue_1; // @[StoreQueue.scala 141:51:@820.4]
  assign _T_1873 = io_loadAddressDone_1 & _T_1872; // @[StoreQueue.scala 141:36:@821.4]
  assign noConflicts_1 = _T_1868 | _T_1873; // @[StoreQueue.scala 140:95:@822.4]
  assign _T_1876 = entriesToCheck_2 == 1'h0; // @[StoreQueue.scala 140:34:@824.4]
  assign _T_1877 = _T_1876 | io_loadDataDone_2; // @[StoreQueue.scala 140:64:@825.4]
  assign _T_1881 = _GEN_263 != io_loadAddressQueue_2; // @[StoreQueue.scala 141:51:@826.4]
  assign _T_1882 = io_loadAddressDone_2 & _T_1881; // @[StoreQueue.scala 141:36:@827.4]
  assign noConflicts_2 = _T_1877 | _T_1882; // @[StoreQueue.scala 140:95:@828.4]
  assign _T_1885 = entriesToCheck_3 == 1'h0; // @[StoreQueue.scala 140:34:@830.4]
  assign _T_1886 = _T_1885 | io_loadDataDone_3; // @[StoreQueue.scala 140:64:@831.4]
  assign _T_1890 = _GEN_263 != io_loadAddressQueue_3; // @[StoreQueue.scala 141:51:@832.4]
  assign _T_1891 = io_loadAddressDone_3 & _T_1890; // @[StoreQueue.scala 141:36:@833.4]
  assign noConflicts_3 = _T_1886 | _T_1891; // @[StoreQueue.scala 140:95:@834.4]
  assign _T_1894 = entriesToCheck_4 == 1'h0; // @[StoreQueue.scala 140:34:@836.4]
  assign _T_1895 = _T_1894 | io_loadDataDone_4; // @[StoreQueue.scala 140:64:@837.4]
  assign _T_1899 = _GEN_263 != io_loadAddressQueue_4; // @[StoreQueue.scala 141:51:@838.4]
  assign _T_1900 = io_loadAddressDone_4 & _T_1899; // @[StoreQueue.scala 141:36:@839.4]
  assign noConflicts_4 = _T_1895 | _T_1900; // @[StoreQueue.scala 140:95:@840.4]
  assign _T_1903 = entriesToCheck_5 == 1'h0; // @[StoreQueue.scala 140:34:@842.4]
  assign _T_1904 = _T_1903 | io_loadDataDone_5; // @[StoreQueue.scala 140:64:@843.4]
  assign _T_1908 = _GEN_263 != io_loadAddressQueue_5; // @[StoreQueue.scala 141:51:@844.4]
  assign _T_1909 = io_loadAddressDone_5 & _T_1908; // @[StoreQueue.scala 141:36:@845.4]
  assign noConflicts_5 = _T_1904 | _T_1909; // @[StoreQueue.scala 140:95:@846.4]
  assign _T_1912 = entriesToCheck_6 == 1'h0; // @[StoreQueue.scala 140:34:@848.4]
  assign _T_1913 = _T_1912 | io_loadDataDone_6; // @[StoreQueue.scala 140:64:@849.4]
  assign _T_1917 = _GEN_263 != io_loadAddressQueue_6; // @[StoreQueue.scala 141:51:@850.4]
  assign _T_1918 = io_loadAddressDone_6 & _T_1917; // @[StoreQueue.scala 141:36:@851.4]
  assign noConflicts_6 = _T_1913 | _T_1918; // @[StoreQueue.scala 140:95:@852.4]
  assign _T_1921 = entriesToCheck_7 == 1'h0; // @[StoreQueue.scala 140:34:@854.4]
  assign _T_1922 = _T_1921 | io_loadDataDone_7; // @[StoreQueue.scala 140:64:@855.4]
  assign _T_1926 = _GEN_263 != io_loadAddressQueue_7; // @[StoreQueue.scala 141:51:@856.4]
  assign _T_1927 = io_loadAddressDone_7 & _T_1926; // @[StoreQueue.scala 141:36:@857.4]
  assign noConflicts_7 = _T_1922 | _T_1927; // @[StoreQueue.scala 140:95:@858.4]
  assign _GEN_265 = 3'h1 == head ? addrKnown_1 : addrKnown_0; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_266 = 3'h2 == head ? addrKnown_2 : _GEN_265; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_267 = 3'h3 == head ? addrKnown_3 : _GEN_266; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_268 = 3'h4 == head ? addrKnown_4 : _GEN_267; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_269 = 3'h5 == head ? addrKnown_5 : _GEN_268; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_270 = 3'h6 == head ? addrKnown_6 : _GEN_269; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_271 = 3'h7 == head ? addrKnown_7 : _GEN_270; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_273 = 3'h1 == head ? dataKnown_1 : dataKnown_0; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_274 = 3'h2 == head ? dataKnown_2 : _GEN_273; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_275 = 3'h3 == head ? dataKnown_3 : _GEN_274; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_276 = 3'h4 == head ? dataKnown_4 : _GEN_275; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_277 = 3'h5 == head ? dataKnown_5 : _GEN_276; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_278 = 3'h6 == head ? dataKnown_6 : _GEN_277; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_279 = 3'h7 == head ? dataKnown_7 : _GEN_278; // @[StoreQueue.scala 154:44:@860.4]
  assign _T_1935 = _GEN_271 & _GEN_279; // @[StoreQueue.scala 154:44:@860.4]
  assign _GEN_281 = 3'h1 == head ? storeCompleted_1 : storeCompleted_0; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_282 = 3'h2 == head ? storeCompleted_2 : _GEN_281; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_283 = 3'h3 == head ? storeCompleted_3 : _GEN_282; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_284 = 3'h4 == head ? storeCompleted_4 : _GEN_283; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_285 = 3'h5 == head ? storeCompleted_5 : _GEN_284; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_286 = 3'h6 == head ? storeCompleted_6 : _GEN_285; // @[StoreQueue.scala 154:66:@861.4]
  assign _GEN_287 = 3'h7 == head ? storeCompleted_7 : _GEN_286; // @[StoreQueue.scala 154:66:@861.4]
  assign _T_1940 = _GEN_287 == 1'h0; // @[StoreQueue.scala 154:66:@861.4]
  assign _T_1941 = _T_1935 & _T_1940; // @[StoreQueue.scala 154:63:@862.4]
  assign _T_1944 = noConflicts_0 & noConflicts_1; // @[StoreQueue.scala 154:109:@864.4]
  assign _T_1945 = _T_1944 & noConflicts_2; // @[StoreQueue.scala 154:109:@865.4]
  assign _T_1946 = _T_1945 & noConflicts_3; // @[StoreQueue.scala 154:109:@866.4]
  assign _T_1947 = _T_1946 & noConflicts_4; // @[StoreQueue.scala 154:109:@867.4]
  assign _T_1948 = _T_1947 & noConflicts_5; // @[StoreQueue.scala 154:109:@868.4]
  assign _T_1949 = _T_1948 & noConflicts_6; // @[StoreQueue.scala 154:109:@869.4]
  assign _T_1950 = _T_1949 & noConflicts_7; // @[StoreQueue.scala 154:109:@870.4]
  assign storeRequest = _T_1941 & _T_1950; // @[StoreQueue.scala 154:88:@871.4]
  assign _T_1953 = head == 3'h0; // @[StoreQueue.scala 164:23:@876.6]
  assign _T_1954 = _T_1953 & storeRequest; // @[StoreQueue.scala 164:43:@877.6]
  assign _T_1955 = _T_1954 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@878.6]
  assign _GEN_288 = _T_1955 ? 1'h1 : storeCompleted_0; // @[StoreQueue.scala 164:86:@879.6]
  assign _GEN_289 = initBits_0 ? 1'h0 : _GEN_288; // @[StoreQueue.scala 162:37:@872.4]
  assign _T_1959 = head == 3'h1; // @[StoreQueue.scala 164:23:@886.6]
  assign _T_1960 = _T_1959 & storeRequest; // @[StoreQueue.scala 164:43:@887.6]
  assign _T_1961 = _T_1960 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@888.6]
  assign _GEN_290 = _T_1961 ? 1'h1 : storeCompleted_1; // @[StoreQueue.scala 164:86:@889.6]
  assign _GEN_291 = initBits_1 ? 1'h0 : _GEN_290; // @[StoreQueue.scala 162:37:@882.4]
  assign _T_1965 = head == 3'h2; // @[StoreQueue.scala 164:23:@896.6]
  assign _T_1966 = _T_1965 & storeRequest; // @[StoreQueue.scala 164:43:@897.6]
  assign _T_1967 = _T_1966 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@898.6]
  assign _GEN_292 = _T_1967 ? 1'h1 : storeCompleted_2; // @[StoreQueue.scala 164:86:@899.6]
  assign _GEN_293 = initBits_2 ? 1'h0 : _GEN_292; // @[StoreQueue.scala 162:37:@892.4]
  assign _T_1971 = head == 3'h3; // @[StoreQueue.scala 164:23:@906.6]
  assign _T_1972 = _T_1971 & storeRequest; // @[StoreQueue.scala 164:43:@907.6]
  assign _T_1973 = _T_1972 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@908.6]
  assign _GEN_294 = _T_1973 ? 1'h1 : storeCompleted_3; // @[StoreQueue.scala 164:86:@909.6]
  assign _GEN_295 = initBits_3 ? 1'h0 : _GEN_294; // @[StoreQueue.scala 162:37:@902.4]
  assign _T_1977 = head == 3'h4; // @[StoreQueue.scala 164:23:@916.6]
  assign _T_1978 = _T_1977 & storeRequest; // @[StoreQueue.scala 164:43:@917.6]
  assign _T_1979 = _T_1978 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@918.6]
  assign _GEN_296 = _T_1979 ? 1'h1 : storeCompleted_4; // @[StoreQueue.scala 164:86:@919.6]
  assign _GEN_297 = initBits_4 ? 1'h0 : _GEN_296; // @[StoreQueue.scala 162:37:@912.4]
  assign _T_1983 = head == 3'h5; // @[StoreQueue.scala 164:23:@926.6]
  assign _T_1984 = _T_1983 & storeRequest; // @[StoreQueue.scala 164:43:@927.6]
  assign _T_1985 = _T_1984 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@928.6]
  assign _GEN_298 = _T_1985 ? 1'h1 : storeCompleted_5; // @[StoreQueue.scala 164:86:@929.6]
  assign _GEN_299 = initBits_5 ? 1'h0 : _GEN_298; // @[StoreQueue.scala 162:37:@922.4]
  assign _T_1989 = head == 3'h6; // @[StoreQueue.scala 164:23:@936.6]
  assign _T_1990 = _T_1989 & storeRequest; // @[StoreQueue.scala 164:43:@937.6]
  assign _T_1991 = _T_1990 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@938.6]
  assign _GEN_300 = _T_1991 ? 1'h1 : storeCompleted_6; // @[StoreQueue.scala 164:86:@939.6]
  assign _GEN_301 = initBits_6 ? 1'h0 : _GEN_300; // @[StoreQueue.scala 162:37:@932.4]
  assign _T_1995 = head == 3'h7; // @[StoreQueue.scala 164:23:@946.6]
  assign _T_1996 = _T_1995 & storeRequest; // @[StoreQueue.scala 164:43:@947.6]
  assign _T_1997 = _T_1996 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@948.6]
  assign _GEN_302 = _T_1997 ? 1'h1 : storeCompleted_7; // @[StoreQueue.scala 164:86:@949.6]
  assign _GEN_303 = initBits_7 ? 1'h0 : _GEN_302; // @[StoreQueue.scala 162:37:@942.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[StoreQueue.scala 180:72:@953.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[StoreQueue.scala 180:72:@955.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[StoreQueue.scala 180:72:@957.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[StoreQueue.scala 180:72:@959.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[StoreQueue.scala 180:72:@961.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[StoreQueue.scala 180:72:@963.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[StoreQueue.scala 180:72:@965.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[StoreQueue.scala 180:72:@967.4]
  assign _T_2410 = addrKnown_0 == 1'h0; // @[StoreQueue.scala 192:91:@987.4]
  assign _T_2411 = entriesPorts_0_0 & _T_2410; // @[StoreQueue.scala 192:88:@988.4]
  assign _T_2413 = addrKnown_1 == 1'h0; // @[StoreQueue.scala 192:91:@989.4]
  assign _T_2414 = entriesPorts_0_1 & _T_2413; // @[StoreQueue.scala 192:88:@990.4]
  assign _T_2416 = addrKnown_2 == 1'h0; // @[StoreQueue.scala 192:91:@991.4]
  assign _T_2417 = entriesPorts_0_2 & _T_2416; // @[StoreQueue.scala 192:88:@992.4]
  assign _T_2419 = addrKnown_3 == 1'h0; // @[StoreQueue.scala 192:91:@993.4]
  assign _T_2420 = entriesPorts_0_3 & _T_2419; // @[StoreQueue.scala 192:88:@994.4]
  assign _T_2422 = addrKnown_4 == 1'h0; // @[StoreQueue.scala 192:91:@995.4]
  assign _T_2423 = entriesPorts_0_4 & _T_2422; // @[StoreQueue.scala 192:88:@996.4]
  assign _T_2425 = addrKnown_5 == 1'h0; // @[StoreQueue.scala 192:91:@997.4]
  assign _T_2426 = entriesPorts_0_5 & _T_2425; // @[StoreQueue.scala 192:88:@998.4]
  assign _T_2428 = addrKnown_6 == 1'h0; // @[StoreQueue.scala 192:91:@999.4]
  assign _T_2429 = entriesPorts_0_6 & _T_2428; // @[StoreQueue.scala 192:88:@1000.4]
  assign _T_2431 = addrKnown_7 == 1'h0; // @[StoreQueue.scala 192:91:@1001.4]
  assign _T_2432 = entriesPorts_0_7 & _T_2431; // @[StoreQueue.scala 192:88:@1002.4]
  assign _T_2448 = dataKnown_0 == 1'h0; // @[StoreQueue.scala 193:91:@1012.4]
  assign _T_2449 = entriesPorts_0_0 & _T_2448; // @[StoreQueue.scala 193:88:@1013.4]
  assign _T_2451 = dataKnown_1 == 1'h0; // @[StoreQueue.scala 193:91:@1014.4]
  assign _T_2452 = entriesPorts_0_1 & _T_2451; // @[StoreQueue.scala 193:88:@1015.4]
  assign _T_2454 = dataKnown_2 == 1'h0; // @[StoreQueue.scala 193:91:@1016.4]
  assign _T_2455 = entriesPorts_0_2 & _T_2454; // @[StoreQueue.scala 193:88:@1017.4]
  assign _T_2457 = dataKnown_3 == 1'h0; // @[StoreQueue.scala 193:91:@1018.4]
  assign _T_2458 = entriesPorts_0_3 & _T_2457; // @[StoreQueue.scala 193:88:@1019.4]
  assign _T_2460 = dataKnown_4 == 1'h0; // @[StoreQueue.scala 193:91:@1020.4]
  assign _T_2461 = entriesPorts_0_4 & _T_2460; // @[StoreQueue.scala 193:88:@1021.4]
  assign _T_2463 = dataKnown_5 == 1'h0; // @[StoreQueue.scala 193:91:@1022.4]
  assign _T_2464 = entriesPorts_0_5 & _T_2463; // @[StoreQueue.scala 193:88:@1023.4]
  assign _T_2466 = dataKnown_6 == 1'h0; // @[StoreQueue.scala 193:91:@1024.4]
  assign _T_2467 = entriesPorts_0_6 & _T_2466; // @[StoreQueue.scala 193:88:@1025.4]
  assign _T_2469 = dataKnown_7 == 1'h0; // @[StoreQueue.scala 193:91:@1026.4]
  assign _T_2470 = entriesPorts_0_7 & _T_2469; // @[StoreQueue.scala 193:88:@1027.4]
  assign _T_2487 = 8'h1 << head; // @[OneHot.scala 52:12:@1038.4]
  assign _T_2489 = _T_2487[0]; // @[util.scala 33:60:@1040.4]
  assign _T_2490 = _T_2487[1]; // @[util.scala 33:60:@1041.4]
  assign _T_2491 = _T_2487[2]; // @[util.scala 33:60:@1042.4]
  assign _T_2492 = _T_2487[3]; // @[util.scala 33:60:@1043.4]
  assign _T_2493 = _T_2487[4]; // @[util.scala 33:60:@1044.4]
  assign _T_2494 = _T_2487[5]; // @[util.scala 33:60:@1045.4]
  assign _T_2495 = _T_2487[6]; // @[util.scala 33:60:@1046.4]
  assign _T_2496 = _T_2487[7]; // @[util.scala 33:60:@1047.4]
  assign _T_2521 = _T_2432 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1057.4]
  assign _T_2522 = _T_2429 ? 8'h40 : _T_2521; // @[Mux.scala 31:69:@1058.4]
  assign _T_2523 = _T_2426 ? 8'h20 : _T_2522; // @[Mux.scala 31:69:@1059.4]
  assign _T_2524 = _T_2423 ? 8'h10 : _T_2523; // @[Mux.scala 31:69:@1060.4]
  assign _T_2525 = _T_2420 ? 8'h8 : _T_2524; // @[Mux.scala 31:69:@1061.4]
  assign _T_2526 = _T_2417 ? 8'h4 : _T_2525; // @[Mux.scala 31:69:@1062.4]
  assign _T_2527 = _T_2414 ? 8'h2 : _T_2526; // @[Mux.scala 31:69:@1063.4]
  assign _T_2528 = _T_2411 ? 8'h1 : _T_2527; // @[Mux.scala 31:69:@1064.4]
  assign _T_2529 = _T_2528[0]; // @[OneHot.scala 66:30:@1065.4]
  assign _T_2530 = _T_2528[1]; // @[OneHot.scala 66:30:@1066.4]
  assign _T_2531 = _T_2528[2]; // @[OneHot.scala 66:30:@1067.4]
  assign _T_2532 = _T_2528[3]; // @[OneHot.scala 66:30:@1068.4]
  assign _T_2533 = _T_2528[4]; // @[OneHot.scala 66:30:@1069.4]
  assign _T_2534 = _T_2528[5]; // @[OneHot.scala 66:30:@1070.4]
  assign _T_2535 = _T_2528[6]; // @[OneHot.scala 66:30:@1071.4]
  assign _T_2536 = _T_2528[7]; // @[OneHot.scala 66:30:@1072.4]
  assign _T_2561 = _T_2411 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1082.4]
  assign _T_2562 = _T_2432 ? 8'h40 : _T_2561; // @[Mux.scala 31:69:@1083.4]
  assign _T_2563 = _T_2429 ? 8'h20 : _T_2562; // @[Mux.scala 31:69:@1084.4]
  assign _T_2564 = _T_2426 ? 8'h10 : _T_2563; // @[Mux.scala 31:69:@1085.4]
  assign _T_2565 = _T_2423 ? 8'h8 : _T_2564; // @[Mux.scala 31:69:@1086.4]
  assign _T_2566 = _T_2420 ? 8'h4 : _T_2565; // @[Mux.scala 31:69:@1087.4]
  assign _T_2567 = _T_2417 ? 8'h2 : _T_2566; // @[Mux.scala 31:69:@1088.4]
  assign _T_2568 = _T_2414 ? 8'h1 : _T_2567; // @[Mux.scala 31:69:@1089.4]
  assign _T_2569 = _T_2568[0]; // @[OneHot.scala 66:30:@1090.4]
  assign _T_2570 = _T_2568[1]; // @[OneHot.scala 66:30:@1091.4]
  assign _T_2571 = _T_2568[2]; // @[OneHot.scala 66:30:@1092.4]
  assign _T_2572 = _T_2568[3]; // @[OneHot.scala 66:30:@1093.4]
  assign _T_2573 = _T_2568[4]; // @[OneHot.scala 66:30:@1094.4]
  assign _T_2574 = _T_2568[5]; // @[OneHot.scala 66:30:@1095.4]
  assign _T_2575 = _T_2568[6]; // @[OneHot.scala 66:30:@1096.4]
  assign _T_2576 = _T_2568[7]; // @[OneHot.scala 66:30:@1097.4]
  assign _T_2601 = _T_2414 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1107.4]
  assign _T_2602 = _T_2411 ? 8'h40 : _T_2601; // @[Mux.scala 31:69:@1108.4]
  assign _T_2603 = _T_2432 ? 8'h20 : _T_2602; // @[Mux.scala 31:69:@1109.4]
  assign _T_2604 = _T_2429 ? 8'h10 : _T_2603; // @[Mux.scala 31:69:@1110.4]
  assign _T_2605 = _T_2426 ? 8'h8 : _T_2604; // @[Mux.scala 31:69:@1111.4]
  assign _T_2606 = _T_2423 ? 8'h4 : _T_2605; // @[Mux.scala 31:69:@1112.4]
  assign _T_2607 = _T_2420 ? 8'h2 : _T_2606; // @[Mux.scala 31:69:@1113.4]
  assign _T_2608 = _T_2417 ? 8'h1 : _T_2607; // @[Mux.scala 31:69:@1114.4]
  assign _T_2609 = _T_2608[0]; // @[OneHot.scala 66:30:@1115.4]
  assign _T_2610 = _T_2608[1]; // @[OneHot.scala 66:30:@1116.4]
  assign _T_2611 = _T_2608[2]; // @[OneHot.scala 66:30:@1117.4]
  assign _T_2612 = _T_2608[3]; // @[OneHot.scala 66:30:@1118.4]
  assign _T_2613 = _T_2608[4]; // @[OneHot.scala 66:30:@1119.4]
  assign _T_2614 = _T_2608[5]; // @[OneHot.scala 66:30:@1120.4]
  assign _T_2615 = _T_2608[6]; // @[OneHot.scala 66:30:@1121.4]
  assign _T_2616 = _T_2608[7]; // @[OneHot.scala 66:30:@1122.4]
  assign _T_2641 = _T_2417 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1132.4]
  assign _T_2642 = _T_2414 ? 8'h40 : _T_2641; // @[Mux.scala 31:69:@1133.4]
  assign _T_2643 = _T_2411 ? 8'h20 : _T_2642; // @[Mux.scala 31:69:@1134.4]
  assign _T_2644 = _T_2432 ? 8'h10 : _T_2643; // @[Mux.scala 31:69:@1135.4]
  assign _T_2645 = _T_2429 ? 8'h8 : _T_2644; // @[Mux.scala 31:69:@1136.4]
  assign _T_2646 = _T_2426 ? 8'h4 : _T_2645; // @[Mux.scala 31:69:@1137.4]
  assign _T_2647 = _T_2423 ? 8'h2 : _T_2646; // @[Mux.scala 31:69:@1138.4]
  assign _T_2648 = _T_2420 ? 8'h1 : _T_2647; // @[Mux.scala 31:69:@1139.4]
  assign _T_2649 = _T_2648[0]; // @[OneHot.scala 66:30:@1140.4]
  assign _T_2650 = _T_2648[1]; // @[OneHot.scala 66:30:@1141.4]
  assign _T_2651 = _T_2648[2]; // @[OneHot.scala 66:30:@1142.4]
  assign _T_2652 = _T_2648[3]; // @[OneHot.scala 66:30:@1143.4]
  assign _T_2653 = _T_2648[4]; // @[OneHot.scala 66:30:@1144.4]
  assign _T_2654 = _T_2648[5]; // @[OneHot.scala 66:30:@1145.4]
  assign _T_2655 = _T_2648[6]; // @[OneHot.scala 66:30:@1146.4]
  assign _T_2656 = _T_2648[7]; // @[OneHot.scala 66:30:@1147.4]
  assign _T_2681 = _T_2420 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1157.4]
  assign _T_2682 = _T_2417 ? 8'h40 : _T_2681; // @[Mux.scala 31:69:@1158.4]
  assign _T_2683 = _T_2414 ? 8'h20 : _T_2682; // @[Mux.scala 31:69:@1159.4]
  assign _T_2684 = _T_2411 ? 8'h10 : _T_2683; // @[Mux.scala 31:69:@1160.4]
  assign _T_2685 = _T_2432 ? 8'h8 : _T_2684; // @[Mux.scala 31:69:@1161.4]
  assign _T_2686 = _T_2429 ? 8'h4 : _T_2685; // @[Mux.scala 31:69:@1162.4]
  assign _T_2687 = _T_2426 ? 8'h2 : _T_2686; // @[Mux.scala 31:69:@1163.4]
  assign _T_2688 = _T_2423 ? 8'h1 : _T_2687; // @[Mux.scala 31:69:@1164.4]
  assign _T_2689 = _T_2688[0]; // @[OneHot.scala 66:30:@1165.4]
  assign _T_2690 = _T_2688[1]; // @[OneHot.scala 66:30:@1166.4]
  assign _T_2691 = _T_2688[2]; // @[OneHot.scala 66:30:@1167.4]
  assign _T_2692 = _T_2688[3]; // @[OneHot.scala 66:30:@1168.4]
  assign _T_2693 = _T_2688[4]; // @[OneHot.scala 66:30:@1169.4]
  assign _T_2694 = _T_2688[5]; // @[OneHot.scala 66:30:@1170.4]
  assign _T_2695 = _T_2688[6]; // @[OneHot.scala 66:30:@1171.4]
  assign _T_2696 = _T_2688[7]; // @[OneHot.scala 66:30:@1172.4]
  assign _T_2721 = _T_2423 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1182.4]
  assign _T_2722 = _T_2420 ? 8'h40 : _T_2721; // @[Mux.scala 31:69:@1183.4]
  assign _T_2723 = _T_2417 ? 8'h20 : _T_2722; // @[Mux.scala 31:69:@1184.4]
  assign _T_2724 = _T_2414 ? 8'h10 : _T_2723; // @[Mux.scala 31:69:@1185.4]
  assign _T_2725 = _T_2411 ? 8'h8 : _T_2724; // @[Mux.scala 31:69:@1186.4]
  assign _T_2726 = _T_2432 ? 8'h4 : _T_2725; // @[Mux.scala 31:69:@1187.4]
  assign _T_2727 = _T_2429 ? 8'h2 : _T_2726; // @[Mux.scala 31:69:@1188.4]
  assign _T_2728 = _T_2426 ? 8'h1 : _T_2727; // @[Mux.scala 31:69:@1189.4]
  assign _T_2729 = _T_2728[0]; // @[OneHot.scala 66:30:@1190.4]
  assign _T_2730 = _T_2728[1]; // @[OneHot.scala 66:30:@1191.4]
  assign _T_2731 = _T_2728[2]; // @[OneHot.scala 66:30:@1192.4]
  assign _T_2732 = _T_2728[3]; // @[OneHot.scala 66:30:@1193.4]
  assign _T_2733 = _T_2728[4]; // @[OneHot.scala 66:30:@1194.4]
  assign _T_2734 = _T_2728[5]; // @[OneHot.scala 66:30:@1195.4]
  assign _T_2735 = _T_2728[6]; // @[OneHot.scala 66:30:@1196.4]
  assign _T_2736 = _T_2728[7]; // @[OneHot.scala 66:30:@1197.4]
  assign _T_2761 = _T_2426 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1207.4]
  assign _T_2762 = _T_2423 ? 8'h40 : _T_2761; // @[Mux.scala 31:69:@1208.4]
  assign _T_2763 = _T_2420 ? 8'h20 : _T_2762; // @[Mux.scala 31:69:@1209.4]
  assign _T_2764 = _T_2417 ? 8'h10 : _T_2763; // @[Mux.scala 31:69:@1210.4]
  assign _T_2765 = _T_2414 ? 8'h8 : _T_2764; // @[Mux.scala 31:69:@1211.4]
  assign _T_2766 = _T_2411 ? 8'h4 : _T_2765; // @[Mux.scala 31:69:@1212.4]
  assign _T_2767 = _T_2432 ? 8'h2 : _T_2766; // @[Mux.scala 31:69:@1213.4]
  assign _T_2768 = _T_2429 ? 8'h1 : _T_2767; // @[Mux.scala 31:69:@1214.4]
  assign _T_2769 = _T_2768[0]; // @[OneHot.scala 66:30:@1215.4]
  assign _T_2770 = _T_2768[1]; // @[OneHot.scala 66:30:@1216.4]
  assign _T_2771 = _T_2768[2]; // @[OneHot.scala 66:30:@1217.4]
  assign _T_2772 = _T_2768[3]; // @[OneHot.scala 66:30:@1218.4]
  assign _T_2773 = _T_2768[4]; // @[OneHot.scala 66:30:@1219.4]
  assign _T_2774 = _T_2768[5]; // @[OneHot.scala 66:30:@1220.4]
  assign _T_2775 = _T_2768[6]; // @[OneHot.scala 66:30:@1221.4]
  assign _T_2776 = _T_2768[7]; // @[OneHot.scala 66:30:@1222.4]
  assign _T_2801 = _T_2429 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1232.4]
  assign _T_2802 = _T_2426 ? 8'h40 : _T_2801; // @[Mux.scala 31:69:@1233.4]
  assign _T_2803 = _T_2423 ? 8'h20 : _T_2802; // @[Mux.scala 31:69:@1234.4]
  assign _T_2804 = _T_2420 ? 8'h10 : _T_2803; // @[Mux.scala 31:69:@1235.4]
  assign _T_2805 = _T_2417 ? 8'h8 : _T_2804; // @[Mux.scala 31:69:@1236.4]
  assign _T_2806 = _T_2414 ? 8'h4 : _T_2805; // @[Mux.scala 31:69:@1237.4]
  assign _T_2807 = _T_2411 ? 8'h2 : _T_2806; // @[Mux.scala 31:69:@1238.4]
  assign _T_2808 = _T_2432 ? 8'h1 : _T_2807; // @[Mux.scala 31:69:@1239.4]
  assign _T_2809 = _T_2808[0]; // @[OneHot.scala 66:30:@1240.4]
  assign _T_2810 = _T_2808[1]; // @[OneHot.scala 66:30:@1241.4]
  assign _T_2811 = _T_2808[2]; // @[OneHot.scala 66:30:@1242.4]
  assign _T_2812 = _T_2808[3]; // @[OneHot.scala 66:30:@1243.4]
  assign _T_2813 = _T_2808[4]; // @[OneHot.scala 66:30:@1244.4]
  assign _T_2814 = _T_2808[5]; // @[OneHot.scala 66:30:@1245.4]
  assign _T_2815 = _T_2808[6]; // @[OneHot.scala 66:30:@1246.4]
  assign _T_2816 = _T_2808[7]; // @[OneHot.scala 66:30:@1247.4]
  assign _T_2857 = {_T_2536,_T_2535,_T_2534,_T_2533,_T_2532,_T_2531,_T_2530,_T_2529}; // @[Mux.scala 19:72:@1263.4]
  assign _T_2859 = _T_2489 ? _T_2857 : 8'h0; // @[Mux.scala 19:72:@1264.4]
  assign _T_2866 = {_T_2575,_T_2574,_T_2573,_T_2572,_T_2571,_T_2570,_T_2569,_T_2576}; // @[Mux.scala 19:72:@1271.4]
  assign _T_2868 = _T_2490 ? _T_2866 : 8'h0; // @[Mux.scala 19:72:@1272.4]
  assign _T_2875 = {_T_2614,_T_2613,_T_2612,_T_2611,_T_2610,_T_2609,_T_2616,_T_2615}; // @[Mux.scala 19:72:@1279.4]
  assign _T_2877 = _T_2491 ? _T_2875 : 8'h0; // @[Mux.scala 19:72:@1280.4]
  assign _T_2884 = {_T_2653,_T_2652,_T_2651,_T_2650,_T_2649,_T_2656,_T_2655,_T_2654}; // @[Mux.scala 19:72:@1287.4]
  assign _T_2886 = _T_2492 ? _T_2884 : 8'h0; // @[Mux.scala 19:72:@1288.4]
  assign _T_2893 = {_T_2692,_T_2691,_T_2690,_T_2689,_T_2696,_T_2695,_T_2694,_T_2693}; // @[Mux.scala 19:72:@1295.4]
  assign _T_2895 = _T_2493 ? _T_2893 : 8'h0; // @[Mux.scala 19:72:@1296.4]
  assign _T_2902 = {_T_2731,_T_2730,_T_2729,_T_2736,_T_2735,_T_2734,_T_2733,_T_2732}; // @[Mux.scala 19:72:@1303.4]
  assign _T_2904 = _T_2494 ? _T_2902 : 8'h0; // @[Mux.scala 19:72:@1304.4]
  assign _T_2911 = {_T_2770,_T_2769,_T_2776,_T_2775,_T_2774,_T_2773,_T_2772,_T_2771}; // @[Mux.scala 19:72:@1311.4]
  assign _T_2913 = _T_2495 ? _T_2911 : 8'h0; // @[Mux.scala 19:72:@1312.4]
  assign _T_2920 = {_T_2809,_T_2816,_T_2815,_T_2814,_T_2813,_T_2812,_T_2811,_T_2810}; // @[Mux.scala 19:72:@1319.4]
  assign _T_2922 = _T_2496 ? _T_2920 : 8'h0; // @[Mux.scala 19:72:@1320.4]
  assign _T_2923 = _T_2859 | _T_2868; // @[Mux.scala 19:72:@1321.4]
  assign _T_2924 = _T_2923 | _T_2877; // @[Mux.scala 19:72:@1322.4]
  assign _T_2925 = _T_2924 | _T_2886; // @[Mux.scala 19:72:@1323.4]
  assign _T_2926 = _T_2925 | _T_2895; // @[Mux.scala 19:72:@1324.4]
  assign _T_2927 = _T_2926 | _T_2904; // @[Mux.scala 19:72:@1325.4]
  assign _T_2928 = _T_2927 | _T_2913; // @[Mux.scala 19:72:@1326.4]
  assign _T_2929 = _T_2928 | _T_2922; // @[Mux.scala 19:72:@1327.4]
  assign inputAddrPriorityPorts_0_0 = _T_2929[0]; // @[Mux.scala 19:72:@1331.4]
  assign inputAddrPriorityPorts_0_1 = _T_2929[1]; // @[Mux.scala 19:72:@1333.4]
  assign inputAddrPriorityPorts_0_2 = _T_2929[2]; // @[Mux.scala 19:72:@1335.4]
  assign inputAddrPriorityPorts_0_3 = _T_2929[3]; // @[Mux.scala 19:72:@1337.4]
  assign inputAddrPriorityPorts_0_4 = _T_2929[4]; // @[Mux.scala 19:72:@1339.4]
  assign inputAddrPriorityPorts_0_5 = _T_2929[5]; // @[Mux.scala 19:72:@1341.4]
  assign inputAddrPriorityPorts_0_6 = _T_2929[6]; // @[Mux.scala 19:72:@1343.4]
  assign inputAddrPriorityPorts_0_7 = _T_2929[7]; // @[Mux.scala 19:72:@1345.4]
  assign _T_3043 = _T_2470 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1375.4]
  assign _T_3044 = _T_2467 ? 8'h40 : _T_3043; // @[Mux.scala 31:69:@1376.4]
  assign _T_3045 = _T_2464 ? 8'h20 : _T_3044; // @[Mux.scala 31:69:@1377.4]
  assign _T_3046 = _T_2461 ? 8'h10 : _T_3045; // @[Mux.scala 31:69:@1378.4]
  assign _T_3047 = _T_2458 ? 8'h8 : _T_3046; // @[Mux.scala 31:69:@1379.4]
  assign _T_3048 = _T_2455 ? 8'h4 : _T_3047; // @[Mux.scala 31:69:@1380.4]
  assign _T_3049 = _T_2452 ? 8'h2 : _T_3048; // @[Mux.scala 31:69:@1381.4]
  assign _T_3050 = _T_2449 ? 8'h1 : _T_3049; // @[Mux.scala 31:69:@1382.4]
  assign _T_3051 = _T_3050[0]; // @[OneHot.scala 66:30:@1383.4]
  assign _T_3052 = _T_3050[1]; // @[OneHot.scala 66:30:@1384.4]
  assign _T_3053 = _T_3050[2]; // @[OneHot.scala 66:30:@1385.4]
  assign _T_3054 = _T_3050[3]; // @[OneHot.scala 66:30:@1386.4]
  assign _T_3055 = _T_3050[4]; // @[OneHot.scala 66:30:@1387.4]
  assign _T_3056 = _T_3050[5]; // @[OneHot.scala 66:30:@1388.4]
  assign _T_3057 = _T_3050[6]; // @[OneHot.scala 66:30:@1389.4]
  assign _T_3058 = _T_3050[7]; // @[OneHot.scala 66:30:@1390.4]
  assign _T_3083 = _T_2449 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1400.4]
  assign _T_3084 = _T_2470 ? 8'h40 : _T_3083; // @[Mux.scala 31:69:@1401.4]
  assign _T_3085 = _T_2467 ? 8'h20 : _T_3084; // @[Mux.scala 31:69:@1402.4]
  assign _T_3086 = _T_2464 ? 8'h10 : _T_3085; // @[Mux.scala 31:69:@1403.4]
  assign _T_3087 = _T_2461 ? 8'h8 : _T_3086; // @[Mux.scala 31:69:@1404.4]
  assign _T_3088 = _T_2458 ? 8'h4 : _T_3087; // @[Mux.scala 31:69:@1405.4]
  assign _T_3089 = _T_2455 ? 8'h2 : _T_3088; // @[Mux.scala 31:69:@1406.4]
  assign _T_3090 = _T_2452 ? 8'h1 : _T_3089; // @[Mux.scala 31:69:@1407.4]
  assign _T_3091 = _T_3090[0]; // @[OneHot.scala 66:30:@1408.4]
  assign _T_3092 = _T_3090[1]; // @[OneHot.scala 66:30:@1409.4]
  assign _T_3093 = _T_3090[2]; // @[OneHot.scala 66:30:@1410.4]
  assign _T_3094 = _T_3090[3]; // @[OneHot.scala 66:30:@1411.4]
  assign _T_3095 = _T_3090[4]; // @[OneHot.scala 66:30:@1412.4]
  assign _T_3096 = _T_3090[5]; // @[OneHot.scala 66:30:@1413.4]
  assign _T_3097 = _T_3090[6]; // @[OneHot.scala 66:30:@1414.4]
  assign _T_3098 = _T_3090[7]; // @[OneHot.scala 66:30:@1415.4]
  assign _T_3123 = _T_2452 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1425.4]
  assign _T_3124 = _T_2449 ? 8'h40 : _T_3123; // @[Mux.scala 31:69:@1426.4]
  assign _T_3125 = _T_2470 ? 8'h20 : _T_3124; // @[Mux.scala 31:69:@1427.4]
  assign _T_3126 = _T_2467 ? 8'h10 : _T_3125; // @[Mux.scala 31:69:@1428.4]
  assign _T_3127 = _T_2464 ? 8'h8 : _T_3126; // @[Mux.scala 31:69:@1429.4]
  assign _T_3128 = _T_2461 ? 8'h4 : _T_3127; // @[Mux.scala 31:69:@1430.4]
  assign _T_3129 = _T_2458 ? 8'h2 : _T_3128; // @[Mux.scala 31:69:@1431.4]
  assign _T_3130 = _T_2455 ? 8'h1 : _T_3129; // @[Mux.scala 31:69:@1432.4]
  assign _T_3131 = _T_3130[0]; // @[OneHot.scala 66:30:@1433.4]
  assign _T_3132 = _T_3130[1]; // @[OneHot.scala 66:30:@1434.4]
  assign _T_3133 = _T_3130[2]; // @[OneHot.scala 66:30:@1435.4]
  assign _T_3134 = _T_3130[3]; // @[OneHot.scala 66:30:@1436.4]
  assign _T_3135 = _T_3130[4]; // @[OneHot.scala 66:30:@1437.4]
  assign _T_3136 = _T_3130[5]; // @[OneHot.scala 66:30:@1438.4]
  assign _T_3137 = _T_3130[6]; // @[OneHot.scala 66:30:@1439.4]
  assign _T_3138 = _T_3130[7]; // @[OneHot.scala 66:30:@1440.4]
  assign _T_3163 = _T_2455 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1450.4]
  assign _T_3164 = _T_2452 ? 8'h40 : _T_3163; // @[Mux.scala 31:69:@1451.4]
  assign _T_3165 = _T_2449 ? 8'h20 : _T_3164; // @[Mux.scala 31:69:@1452.4]
  assign _T_3166 = _T_2470 ? 8'h10 : _T_3165; // @[Mux.scala 31:69:@1453.4]
  assign _T_3167 = _T_2467 ? 8'h8 : _T_3166; // @[Mux.scala 31:69:@1454.4]
  assign _T_3168 = _T_2464 ? 8'h4 : _T_3167; // @[Mux.scala 31:69:@1455.4]
  assign _T_3169 = _T_2461 ? 8'h2 : _T_3168; // @[Mux.scala 31:69:@1456.4]
  assign _T_3170 = _T_2458 ? 8'h1 : _T_3169; // @[Mux.scala 31:69:@1457.4]
  assign _T_3171 = _T_3170[0]; // @[OneHot.scala 66:30:@1458.4]
  assign _T_3172 = _T_3170[1]; // @[OneHot.scala 66:30:@1459.4]
  assign _T_3173 = _T_3170[2]; // @[OneHot.scala 66:30:@1460.4]
  assign _T_3174 = _T_3170[3]; // @[OneHot.scala 66:30:@1461.4]
  assign _T_3175 = _T_3170[4]; // @[OneHot.scala 66:30:@1462.4]
  assign _T_3176 = _T_3170[5]; // @[OneHot.scala 66:30:@1463.4]
  assign _T_3177 = _T_3170[6]; // @[OneHot.scala 66:30:@1464.4]
  assign _T_3178 = _T_3170[7]; // @[OneHot.scala 66:30:@1465.4]
  assign _T_3203 = _T_2458 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1475.4]
  assign _T_3204 = _T_2455 ? 8'h40 : _T_3203; // @[Mux.scala 31:69:@1476.4]
  assign _T_3205 = _T_2452 ? 8'h20 : _T_3204; // @[Mux.scala 31:69:@1477.4]
  assign _T_3206 = _T_2449 ? 8'h10 : _T_3205; // @[Mux.scala 31:69:@1478.4]
  assign _T_3207 = _T_2470 ? 8'h8 : _T_3206; // @[Mux.scala 31:69:@1479.4]
  assign _T_3208 = _T_2467 ? 8'h4 : _T_3207; // @[Mux.scala 31:69:@1480.4]
  assign _T_3209 = _T_2464 ? 8'h2 : _T_3208; // @[Mux.scala 31:69:@1481.4]
  assign _T_3210 = _T_2461 ? 8'h1 : _T_3209; // @[Mux.scala 31:69:@1482.4]
  assign _T_3211 = _T_3210[0]; // @[OneHot.scala 66:30:@1483.4]
  assign _T_3212 = _T_3210[1]; // @[OneHot.scala 66:30:@1484.4]
  assign _T_3213 = _T_3210[2]; // @[OneHot.scala 66:30:@1485.4]
  assign _T_3214 = _T_3210[3]; // @[OneHot.scala 66:30:@1486.4]
  assign _T_3215 = _T_3210[4]; // @[OneHot.scala 66:30:@1487.4]
  assign _T_3216 = _T_3210[5]; // @[OneHot.scala 66:30:@1488.4]
  assign _T_3217 = _T_3210[6]; // @[OneHot.scala 66:30:@1489.4]
  assign _T_3218 = _T_3210[7]; // @[OneHot.scala 66:30:@1490.4]
  assign _T_3243 = _T_2461 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1500.4]
  assign _T_3244 = _T_2458 ? 8'h40 : _T_3243; // @[Mux.scala 31:69:@1501.4]
  assign _T_3245 = _T_2455 ? 8'h20 : _T_3244; // @[Mux.scala 31:69:@1502.4]
  assign _T_3246 = _T_2452 ? 8'h10 : _T_3245; // @[Mux.scala 31:69:@1503.4]
  assign _T_3247 = _T_2449 ? 8'h8 : _T_3246; // @[Mux.scala 31:69:@1504.4]
  assign _T_3248 = _T_2470 ? 8'h4 : _T_3247; // @[Mux.scala 31:69:@1505.4]
  assign _T_3249 = _T_2467 ? 8'h2 : _T_3248; // @[Mux.scala 31:69:@1506.4]
  assign _T_3250 = _T_2464 ? 8'h1 : _T_3249; // @[Mux.scala 31:69:@1507.4]
  assign _T_3251 = _T_3250[0]; // @[OneHot.scala 66:30:@1508.4]
  assign _T_3252 = _T_3250[1]; // @[OneHot.scala 66:30:@1509.4]
  assign _T_3253 = _T_3250[2]; // @[OneHot.scala 66:30:@1510.4]
  assign _T_3254 = _T_3250[3]; // @[OneHot.scala 66:30:@1511.4]
  assign _T_3255 = _T_3250[4]; // @[OneHot.scala 66:30:@1512.4]
  assign _T_3256 = _T_3250[5]; // @[OneHot.scala 66:30:@1513.4]
  assign _T_3257 = _T_3250[6]; // @[OneHot.scala 66:30:@1514.4]
  assign _T_3258 = _T_3250[7]; // @[OneHot.scala 66:30:@1515.4]
  assign _T_3283 = _T_2464 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1525.4]
  assign _T_3284 = _T_2461 ? 8'h40 : _T_3283; // @[Mux.scala 31:69:@1526.4]
  assign _T_3285 = _T_2458 ? 8'h20 : _T_3284; // @[Mux.scala 31:69:@1527.4]
  assign _T_3286 = _T_2455 ? 8'h10 : _T_3285; // @[Mux.scala 31:69:@1528.4]
  assign _T_3287 = _T_2452 ? 8'h8 : _T_3286; // @[Mux.scala 31:69:@1529.4]
  assign _T_3288 = _T_2449 ? 8'h4 : _T_3287; // @[Mux.scala 31:69:@1530.4]
  assign _T_3289 = _T_2470 ? 8'h2 : _T_3288; // @[Mux.scala 31:69:@1531.4]
  assign _T_3290 = _T_2467 ? 8'h1 : _T_3289; // @[Mux.scala 31:69:@1532.4]
  assign _T_3291 = _T_3290[0]; // @[OneHot.scala 66:30:@1533.4]
  assign _T_3292 = _T_3290[1]; // @[OneHot.scala 66:30:@1534.4]
  assign _T_3293 = _T_3290[2]; // @[OneHot.scala 66:30:@1535.4]
  assign _T_3294 = _T_3290[3]; // @[OneHot.scala 66:30:@1536.4]
  assign _T_3295 = _T_3290[4]; // @[OneHot.scala 66:30:@1537.4]
  assign _T_3296 = _T_3290[5]; // @[OneHot.scala 66:30:@1538.4]
  assign _T_3297 = _T_3290[6]; // @[OneHot.scala 66:30:@1539.4]
  assign _T_3298 = _T_3290[7]; // @[OneHot.scala 66:30:@1540.4]
  assign _T_3323 = _T_2467 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1550.4]
  assign _T_3324 = _T_2464 ? 8'h40 : _T_3323; // @[Mux.scala 31:69:@1551.4]
  assign _T_3325 = _T_2461 ? 8'h20 : _T_3324; // @[Mux.scala 31:69:@1552.4]
  assign _T_3326 = _T_2458 ? 8'h10 : _T_3325; // @[Mux.scala 31:69:@1553.4]
  assign _T_3327 = _T_2455 ? 8'h8 : _T_3326; // @[Mux.scala 31:69:@1554.4]
  assign _T_3328 = _T_2452 ? 8'h4 : _T_3327; // @[Mux.scala 31:69:@1555.4]
  assign _T_3329 = _T_2449 ? 8'h2 : _T_3328; // @[Mux.scala 31:69:@1556.4]
  assign _T_3330 = _T_2470 ? 8'h1 : _T_3329; // @[Mux.scala 31:69:@1557.4]
  assign _T_3331 = _T_3330[0]; // @[OneHot.scala 66:30:@1558.4]
  assign _T_3332 = _T_3330[1]; // @[OneHot.scala 66:30:@1559.4]
  assign _T_3333 = _T_3330[2]; // @[OneHot.scala 66:30:@1560.4]
  assign _T_3334 = _T_3330[3]; // @[OneHot.scala 66:30:@1561.4]
  assign _T_3335 = _T_3330[4]; // @[OneHot.scala 66:30:@1562.4]
  assign _T_3336 = _T_3330[5]; // @[OneHot.scala 66:30:@1563.4]
  assign _T_3337 = _T_3330[6]; // @[OneHot.scala 66:30:@1564.4]
  assign _T_3338 = _T_3330[7]; // @[OneHot.scala 66:30:@1565.4]
  assign _T_3379 = {_T_3058,_T_3057,_T_3056,_T_3055,_T_3054,_T_3053,_T_3052,_T_3051}; // @[Mux.scala 19:72:@1581.4]
  assign _T_3381 = _T_2489 ? _T_3379 : 8'h0; // @[Mux.scala 19:72:@1582.4]
  assign _T_3388 = {_T_3097,_T_3096,_T_3095,_T_3094,_T_3093,_T_3092,_T_3091,_T_3098}; // @[Mux.scala 19:72:@1589.4]
  assign _T_3390 = _T_2490 ? _T_3388 : 8'h0; // @[Mux.scala 19:72:@1590.4]
  assign _T_3397 = {_T_3136,_T_3135,_T_3134,_T_3133,_T_3132,_T_3131,_T_3138,_T_3137}; // @[Mux.scala 19:72:@1597.4]
  assign _T_3399 = _T_2491 ? _T_3397 : 8'h0; // @[Mux.scala 19:72:@1598.4]
  assign _T_3406 = {_T_3175,_T_3174,_T_3173,_T_3172,_T_3171,_T_3178,_T_3177,_T_3176}; // @[Mux.scala 19:72:@1605.4]
  assign _T_3408 = _T_2492 ? _T_3406 : 8'h0; // @[Mux.scala 19:72:@1606.4]
  assign _T_3415 = {_T_3214,_T_3213,_T_3212,_T_3211,_T_3218,_T_3217,_T_3216,_T_3215}; // @[Mux.scala 19:72:@1613.4]
  assign _T_3417 = _T_2493 ? _T_3415 : 8'h0; // @[Mux.scala 19:72:@1614.4]
  assign _T_3424 = {_T_3253,_T_3252,_T_3251,_T_3258,_T_3257,_T_3256,_T_3255,_T_3254}; // @[Mux.scala 19:72:@1621.4]
  assign _T_3426 = _T_2494 ? _T_3424 : 8'h0; // @[Mux.scala 19:72:@1622.4]
  assign _T_3433 = {_T_3292,_T_3291,_T_3298,_T_3297,_T_3296,_T_3295,_T_3294,_T_3293}; // @[Mux.scala 19:72:@1629.4]
  assign _T_3435 = _T_2495 ? _T_3433 : 8'h0; // @[Mux.scala 19:72:@1630.4]
  assign _T_3442 = {_T_3331,_T_3338,_T_3337,_T_3336,_T_3335,_T_3334,_T_3333,_T_3332}; // @[Mux.scala 19:72:@1637.4]
  assign _T_3444 = _T_2496 ? _T_3442 : 8'h0; // @[Mux.scala 19:72:@1638.4]
  assign _T_3445 = _T_3381 | _T_3390; // @[Mux.scala 19:72:@1639.4]
  assign _T_3446 = _T_3445 | _T_3399; // @[Mux.scala 19:72:@1640.4]
  assign _T_3447 = _T_3446 | _T_3408; // @[Mux.scala 19:72:@1641.4]
  assign _T_3448 = _T_3447 | _T_3417; // @[Mux.scala 19:72:@1642.4]
  assign _T_3449 = _T_3448 | _T_3426; // @[Mux.scala 19:72:@1643.4]
  assign _T_3450 = _T_3449 | _T_3435; // @[Mux.scala 19:72:@1644.4]
  assign _T_3451 = _T_3450 | _T_3444; // @[Mux.scala 19:72:@1645.4]
  assign inputDataPriorityPorts_0_0 = _T_3451[0]; // @[Mux.scala 19:72:@1649.4]
  assign inputDataPriorityPorts_0_1 = _T_3451[1]; // @[Mux.scala 19:72:@1651.4]
  assign inputDataPriorityPorts_0_2 = _T_3451[2]; // @[Mux.scala 19:72:@1653.4]
  assign inputDataPriorityPorts_0_3 = _T_3451[3]; // @[Mux.scala 19:72:@1655.4]
  assign inputDataPriorityPorts_0_4 = _T_3451[4]; // @[Mux.scala 19:72:@1657.4]
  assign inputDataPriorityPorts_0_5 = _T_3451[5]; // @[Mux.scala 19:72:@1659.4]
  assign inputDataPriorityPorts_0_6 = _T_3451[6]; // @[Mux.scala 19:72:@1661.4]
  assign inputDataPriorityPorts_0_7 = _T_3451[7]; // @[Mux.scala 19:72:@1663.4]
  assign _T_3531 = portQ_0 & _T_2410; // @[StoreQueue.scala 192:88:@1674.4]
  assign _T_3534 = portQ_1 & _T_2413; // @[StoreQueue.scala 192:88:@1676.4]
  assign _T_3537 = portQ_2 & _T_2416; // @[StoreQueue.scala 192:88:@1678.4]
  assign _T_3540 = portQ_3 & _T_2419; // @[StoreQueue.scala 192:88:@1680.4]
  assign _T_3543 = portQ_4 & _T_2422; // @[StoreQueue.scala 192:88:@1682.4]
  assign _T_3546 = portQ_5 & _T_2425; // @[StoreQueue.scala 192:88:@1684.4]
  assign _T_3549 = portQ_6 & _T_2428; // @[StoreQueue.scala 192:88:@1686.4]
  assign _T_3552 = portQ_7 & _T_2431; // @[StoreQueue.scala 192:88:@1688.4]
  assign _T_3569 = portQ_0 & _T_2448; // @[StoreQueue.scala 193:88:@1699.4]
  assign _T_3572 = portQ_1 & _T_2451; // @[StoreQueue.scala 193:88:@1701.4]
  assign _T_3575 = portQ_2 & _T_2454; // @[StoreQueue.scala 193:88:@1703.4]
  assign _T_3578 = portQ_3 & _T_2457; // @[StoreQueue.scala 193:88:@1705.4]
  assign _T_3581 = portQ_4 & _T_2460; // @[StoreQueue.scala 193:88:@1707.4]
  assign _T_3584 = portQ_5 & _T_2463; // @[StoreQueue.scala 193:88:@1709.4]
  assign _T_3587 = portQ_6 & _T_2466; // @[StoreQueue.scala 193:88:@1711.4]
  assign _T_3590 = portQ_7 & _T_2469; // @[StoreQueue.scala 193:88:@1713.4]
  assign _T_3641 = _T_3552 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1743.4]
  assign _T_3642 = _T_3549 ? 8'h40 : _T_3641; // @[Mux.scala 31:69:@1744.4]
  assign _T_3643 = _T_3546 ? 8'h20 : _T_3642; // @[Mux.scala 31:69:@1745.4]
  assign _T_3644 = _T_3543 ? 8'h10 : _T_3643; // @[Mux.scala 31:69:@1746.4]
  assign _T_3645 = _T_3540 ? 8'h8 : _T_3644; // @[Mux.scala 31:69:@1747.4]
  assign _T_3646 = _T_3537 ? 8'h4 : _T_3645; // @[Mux.scala 31:69:@1748.4]
  assign _T_3647 = _T_3534 ? 8'h2 : _T_3646; // @[Mux.scala 31:69:@1749.4]
  assign _T_3648 = _T_3531 ? 8'h1 : _T_3647; // @[Mux.scala 31:69:@1750.4]
  assign _T_3649 = _T_3648[0]; // @[OneHot.scala 66:30:@1751.4]
  assign _T_3650 = _T_3648[1]; // @[OneHot.scala 66:30:@1752.4]
  assign _T_3651 = _T_3648[2]; // @[OneHot.scala 66:30:@1753.4]
  assign _T_3652 = _T_3648[3]; // @[OneHot.scala 66:30:@1754.4]
  assign _T_3653 = _T_3648[4]; // @[OneHot.scala 66:30:@1755.4]
  assign _T_3654 = _T_3648[5]; // @[OneHot.scala 66:30:@1756.4]
  assign _T_3655 = _T_3648[6]; // @[OneHot.scala 66:30:@1757.4]
  assign _T_3656 = _T_3648[7]; // @[OneHot.scala 66:30:@1758.4]
  assign _T_3681 = _T_3531 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1768.4]
  assign _T_3682 = _T_3552 ? 8'h40 : _T_3681; // @[Mux.scala 31:69:@1769.4]
  assign _T_3683 = _T_3549 ? 8'h20 : _T_3682; // @[Mux.scala 31:69:@1770.4]
  assign _T_3684 = _T_3546 ? 8'h10 : _T_3683; // @[Mux.scala 31:69:@1771.4]
  assign _T_3685 = _T_3543 ? 8'h8 : _T_3684; // @[Mux.scala 31:69:@1772.4]
  assign _T_3686 = _T_3540 ? 8'h4 : _T_3685; // @[Mux.scala 31:69:@1773.4]
  assign _T_3687 = _T_3537 ? 8'h2 : _T_3686; // @[Mux.scala 31:69:@1774.4]
  assign _T_3688 = _T_3534 ? 8'h1 : _T_3687; // @[Mux.scala 31:69:@1775.4]
  assign _T_3689 = _T_3688[0]; // @[OneHot.scala 66:30:@1776.4]
  assign _T_3690 = _T_3688[1]; // @[OneHot.scala 66:30:@1777.4]
  assign _T_3691 = _T_3688[2]; // @[OneHot.scala 66:30:@1778.4]
  assign _T_3692 = _T_3688[3]; // @[OneHot.scala 66:30:@1779.4]
  assign _T_3693 = _T_3688[4]; // @[OneHot.scala 66:30:@1780.4]
  assign _T_3694 = _T_3688[5]; // @[OneHot.scala 66:30:@1781.4]
  assign _T_3695 = _T_3688[6]; // @[OneHot.scala 66:30:@1782.4]
  assign _T_3696 = _T_3688[7]; // @[OneHot.scala 66:30:@1783.4]
  assign _T_3721 = _T_3534 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1793.4]
  assign _T_3722 = _T_3531 ? 8'h40 : _T_3721; // @[Mux.scala 31:69:@1794.4]
  assign _T_3723 = _T_3552 ? 8'h20 : _T_3722; // @[Mux.scala 31:69:@1795.4]
  assign _T_3724 = _T_3549 ? 8'h10 : _T_3723; // @[Mux.scala 31:69:@1796.4]
  assign _T_3725 = _T_3546 ? 8'h8 : _T_3724; // @[Mux.scala 31:69:@1797.4]
  assign _T_3726 = _T_3543 ? 8'h4 : _T_3725; // @[Mux.scala 31:69:@1798.4]
  assign _T_3727 = _T_3540 ? 8'h2 : _T_3726; // @[Mux.scala 31:69:@1799.4]
  assign _T_3728 = _T_3537 ? 8'h1 : _T_3727; // @[Mux.scala 31:69:@1800.4]
  assign _T_3729 = _T_3728[0]; // @[OneHot.scala 66:30:@1801.4]
  assign _T_3730 = _T_3728[1]; // @[OneHot.scala 66:30:@1802.4]
  assign _T_3731 = _T_3728[2]; // @[OneHot.scala 66:30:@1803.4]
  assign _T_3732 = _T_3728[3]; // @[OneHot.scala 66:30:@1804.4]
  assign _T_3733 = _T_3728[4]; // @[OneHot.scala 66:30:@1805.4]
  assign _T_3734 = _T_3728[5]; // @[OneHot.scala 66:30:@1806.4]
  assign _T_3735 = _T_3728[6]; // @[OneHot.scala 66:30:@1807.4]
  assign _T_3736 = _T_3728[7]; // @[OneHot.scala 66:30:@1808.4]
  assign _T_3761 = _T_3537 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1818.4]
  assign _T_3762 = _T_3534 ? 8'h40 : _T_3761; // @[Mux.scala 31:69:@1819.4]
  assign _T_3763 = _T_3531 ? 8'h20 : _T_3762; // @[Mux.scala 31:69:@1820.4]
  assign _T_3764 = _T_3552 ? 8'h10 : _T_3763; // @[Mux.scala 31:69:@1821.4]
  assign _T_3765 = _T_3549 ? 8'h8 : _T_3764; // @[Mux.scala 31:69:@1822.4]
  assign _T_3766 = _T_3546 ? 8'h4 : _T_3765; // @[Mux.scala 31:69:@1823.4]
  assign _T_3767 = _T_3543 ? 8'h2 : _T_3766; // @[Mux.scala 31:69:@1824.4]
  assign _T_3768 = _T_3540 ? 8'h1 : _T_3767; // @[Mux.scala 31:69:@1825.4]
  assign _T_3769 = _T_3768[0]; // @[OneHot.scala 66:30:@1826.4]
  assign _T_3770 = _T_3768[1]; // @[OneHot.scala 66:30:@1827.4]
  assign _T_3771 = _T_3768[2]; // @[OneHot.scala 66:30:@1828.4]
  assign _T_3772 = _T_3768[3]; // @[OneHot.scala 66:30:@1829.4]
  assign _T_3773 = _T_3768[4]; // @[OneHot.scala 66:30:@1830.4]
  assign _T_3774 = _T_3768[5]; // @[OneHot.scala 66:30:@1831.4]
  assign _T_3775 = _T_3768[6]; // @[OneHot.scala 66:30:@1832.4]
  assign _T_3776 = _T_3768[7]; // @[OneHot.scala 66:30:@1833.4]
  assign _T_3801 = _T_3540 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1843.4]
  assign _T_3802 = _T_3537 ? 8'h40 : _T_3801; // @[Mux.scala 31:69:@1844.4]
  assign _T_3803 = _T_3534 ? 8'h20 : _T_3802; // @[Mux.scala 31:69:@1845.4]
  assign _T_3804 = _T_3531 ? 8'h10 : _T_3803; // @[Mux.scala 31:69:@1846.4]
  assign _T_3805 = _T_3552 ? 8'h8 : _T_3804; // @[Mux.scala 31:69:@1847.4]
  assign _T_3806 = _T_3549 ? 8'h4 : _T_3805; // @[Mux.scala 31:69:@1848.4]
  assign _T_3807 = _T_3546 ? 8'h2 : _T_3806; // @[Mux.scala 31:69:@1849.4]
  assign _T_3808 = _T_3543 ? 8'h1 : _T_3807; // @[Mux.scala 31:69:@1850.4]
  assign _T_3809 = _T_3808[0]; // @[OneHot.scala 66:30:@1851.4]
  assign _T_3810 = _T_3808[1]; // @[OneHot.scala 66:30:@1852.4]
  assign _T_3811 = _T_3808[2]; // @[OneHot.scala 66:30:@1853.4]
  assign _T_3812 = _T_3808[3]; // @[OneHot.scala 66:30:@1854.4]
  assign _T_3813 = _T_3808[4]; // @[OneHot.scala 66:30:@1855.4]
  assign _T_3814 = _T_3808[5]; // @[OneHot.scala 66:30:@1856.4]
  assign _T_3815 = _T_3808[6]; // @[OneHot.scala 66:30:@1857.4]
  assign _T_3816 = _T_3808[7]; // @[OneHot.scala 66:30:@1858.4]
  assign _T_3841 = _T_3543 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1868.4]
  assign _T_3842 = _T_3540 ? 8'h40 : _T_3841; // @[Mux.scala 31:69:@1869.4]
  assign _T_3843 = _T_3537 ? 8'h20 : _T_3842; // @[Mux.scala 31:69:@1870.4]
  assign _T_3844 = _T_3534 ? 8'h10 : _T_3843; // @[Mux.scala 31:69:@1871.4]
  assign _T_3845 = _T_3531 ? 8'h8 : _T_3844; // @[Mux.scala 31:69:@1872.4]
  assign _T_3846 = _T_3552 ? 8'h4 : _T_3845; // @[Mux.scala 31:69:@1873.4]
  assign _T_3847 = _T_3549 ? 8'h2 : _T_3846; // @[Mux.scala 31:69:@1874.4]
  assign _T_3848 = _T_3546 ? 8'h1 : _T_3847; // @[Mux.scala 31:69:@1875.4]
  assign _T_3849 = _T_3848[0]; // @[OneHot.scala 66:30:@1876.4]
  assign _T_3850 = _T_3848[1]; // @[OneHot.scala 66:30:@1877.4]
  assign _T_3851 = _T_3848[2]; // @[OneHot.scala 66:30:@1878.4]
  assign _T_3852 = _T_3848[3]; // @[OneHot.scala 66:30:@1879.4]
  assign _T_3853 = _T_3848[4]; // @[OneHot.scala 66:30:@1880.4]
  assign _T_3854 = _T_3848[5]; // @[OneHot.scala 66:30:@1881.4]
  assign _T_3855 = _T_3848[6]; // @[OneHot.scala 66:30:@1882.4]
  assign _T_3856 = _T_3848[7]; // @[OneHot.scala 66:30:@1883.4]
  assign _T_3881 = _T_3546 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1893.4]
  assign _T_3882 = _T_3543 ? 8'h40 : _T_3881; // @[Mux.scala 31:69:@1894.4]
  assign _T_3883 = _T_3540 ? 8'h20 : _T_3882; // @[Mux.scala 31:69:@1895.4]
  assign _T_3884 = _T_3537 ? 8'h10 : _T_3883; // @[Mux.scala 31:69:@1896.4]
  assign _T_3885 = _T_3534 ? 8'h8 : _T_3884; // @[Mux.scala 31:69:@1897.4]
  assign _T_3886 = _T_3531 ? 8'h4 : _T_3885; // @[Mux.scala 31:69:@1898.4]
  assign _T_3887 = _T_3552 ? 8'h2 : _T_3886; // @[Mux.scala 31:69:@1899.4]
  assign _T_3888 = _T_3549 ? 8'h1 : _T_3887; // @[Mux.scala 31:69:@1900.4]
  assign _T_3889 = _T_3888[0]; // @[OneHot.scala 66:30:@1901.4]
  assign _T_3890 = _T_3888[1]; // @[OneHot.scala 66:30:@1902.4]
  assign _T_3891 = _T_3888[2]; // @[OneHot.scala 66:30:@1903.4]
  assign _T_3892 = _T_3888[3]; // @[OneHot.scala 66:30:@1904.4]
  assign _T_3893 = _T_3888[4]; // @[OneHot.scala 66:30:@1905.4]
  assign _T_3894 = _T_3888[5]; // @[OneHot.scala 66:30:@1906.4]
  assign _T_3895 = _T_3888[6]; // @[OneHot.scala 66:30:@1907.4]
  assign _T_3896 = _T_3888[7]; // @[OneHot.scala 66:30:@1908.4]
  assign _T_3921 = _T_3549 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@1918.4]
  assign _T_3922 = _T_3546 ? 8'h40 : _T_3921; // @[Mux.scala 31:69:@1919.4]
  assign _T_3923 = _T_3543 ? 8'h20 : _T_3922; // @[Mux.scala 31:69:@1920.4]
  assign _T_3924 = _T_3540 ? 8'h10 : _T_3923; // @[Mux.scala 31:69:@1921.4]
  assign _T_3925 = _T_3537 ? 8'h8 : _T_3924; // @[Mux.scala 31:69:@1922.4]
  assign _T_3926 = _T_3534 ? 8'h4 : _T_3925; // @[Mux.scala 31:69:@1923.4]
  assign _T_3927 = _T_3531 ? 8'h2 : _T_3926; // @[Mux.scala 31:69:@1924.4]
  assign _T_3928 = _T_3552 ? 8'h1 : _T_3927; // @[Mux.scala 31:69:@1925.4]
  assign _T_3929 = _T_3928[0]; // @[OneHot.scala 66:30:@1926.4]
  assign _T_3930 = _T_3928[1]; // @[OneHot.scala 66:30:@1927.4]
  assign _T_3931 = _T_3928[2]; // @[OneHot.scala 66:30:@1928.4]
  assign _T_3932 = _T_3928[3]; // @[OneHot.scala 66:30:@1929.4]
  assign _T_3933 = _T_3928[4]; // @[OneHot.scala 66:30:@1930.4]
  assign _T_3934 = _T_3928[5]; // @[OneHot.scala 66:30:@1931.4]
  assign _T_3935 = _T_3928[6]; // @[OneHot.scala 66:30:@1932.4]
  assign _T_3936 = _T_3928[7]; // @[OneHot.scala 66:30:@1933.4]
  assign _T_3977 = {_T_3656,_T_3655,_T_3654,_T_3653,_T_3652,_T_3651,_T_3650,_T_3649}; // @[Mux.scala 19:72:@1949.4]
  assign _T_3979 = _T_2489 ? _T_3977 : 8'h0; // @[Mux.scala 19:72:@1950.4]
  assign _T_3986 = {_T_3695,_T_3694,_T_3693,_T_3692,_T_3691,_T_3690,_T_3689,_T_3696}; // @[Mux.scala 19:72:@1957.4]
  assign _T_3988 = _T_2490 ? _T_3986 : 8'h0; // @[Mux.scala 19:72:@1958.4]
  assign _T_3995 = {_T_3734,_T_3733,_T_3732,_T_3731,_T_3730,_T_3729,_T_3736,_T_3735}; // @[Mux.scala 19:72:@1965.4]
  assign _T_3997 = _T_2491 ? _T_3995 : 8'h0; // @[Mux.scala 19:72:@1966.4]
  assign _T_4004 = {_T_3773,_T_3772,_T_3771,_T_3770,_T_3769,_T_3776,_T_3775,_T_3774}; // @[Mux.scala 19:72:@1973.4]
  assign _T_4006 = _T_2492 ? _T_4004 : 8'h0; // @[Mux.scala 19:72:@1974.4]
  assign _T_4013 = {_T_3812,_T_3811,_T_3810,_T_3809,_T_3816,_T_3815,_T_3814,_T_3813}; // @[Mux.scala 19:72:@1981.4]
  assign _T_4015 = _T_2493 ? _T_4013 : 8'h0; // @[Mux.scala 19:72:@1982.4]
  assign _T_4022 = {_T_3851,_T_3850,_T_3849,_T_3856,_T_3855,_T_3854,_T_3853,_T_3852}; // @[Mux.scala 19:72:@1989.4]
  assign _T_4024 = _T_2494 ? _T_4022 : 8'h0; // @[Mux.scala 19:72:@1990.4]
  assign _T_4031 = {_T_3890,_T_3889,_T_3896,_T_3895,_T_3894,_T_3893,_T_3892,_T_3891}; // @[Mux.scala 19:72:@1997.4]
  assign _T_4033 = _T_2495 ? _T_4031 : 8'h0; // @[Mux.scala 19:72:@1998.4]
  assign _T_4040 = {_T_3929,_T_3936,_T_3935,_T_3934,_T_3933,_T_3932,_T_3931,_T_3930}; // @[Mux.scala 19:72:@2005.4]
  assign _T_4042 = _T_2496 ? _T_4040 : 8'h0; // @[Mux.scala 19:72:@2006.4]
  assign _T_4043 = _T_3979 | _T_3988; // @[Mux.scala 19:72:@2007.4]
  assign _T_4044 = _T_4043 | _T_3997; // @[Mux.scala 19:72:@2008.4]
  assign _T_4045 = _T_4044 | _T_4006; // @[Mux.scala 19:72:@2009.4]
  assign _T_4046 = _T_4045 | _T_4015; // @[Mux.scala 19:72:@2010.4]
  assign _T_4047 = _T_4046 | _T_4024; // @[Mux.scala 19:72:@2011.4]
  assign _T_4048 = _T_4047 | _T_4033; // @[Mux.scala 19:72:@2012.4]
  assign _T_4049 = _T_4048 | _T_4042; // @[Mux.scala 19:72:@2013.4]
  assign inputAddrPriorityPorts_1_0 = _T_4049[0]; // @[Mux.scala 19:72:@2017.4]
  assign inputAddrPriorityPorts_1_1 = _T_4049[1]; // @[Mux.scala 19:72:@2019.4]
  assign inputAddrPriorityPorts_1_2 = _T_4049[2]; // @[Mux.scala 19:72:@2021.4]
  assign inputAddrPriorityPorts_1_3 = _T_4049[3]; // @[Mux.scala 19:72:@2023.4]
  assign inputAddrPriorityPorts_1_4 = _T_4049[4]; // @[Mux.scala 19:72:@2025.4]
  assign inputAddrPriorityPorts_1_5 = _T_4049[5]; // @[Mux.scala 19:72:@2027.4]
  assign inputAddrPriorityPorts_1_6 = _T_4049[6]; // @[Mux.scala 19:72:@2029.4]
  assign inputAddrPriorityPorts_1_7 = _T_4049[7]; // @[Mux.scala 19:72:@2031.4]
  assign _T_4163 = _T_3590 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@2061.4]
  assign _T_4164 = _T_3587 ? 8'h40 : _T_4163; // @[Mux.scala 31:69:@2062.4]
  assign _T_4165 = _T_3584 ? 8'h20 : _T_4164; // @[Mux.scala 31:69:@2063.4]
  assign _T_4166 = _T_3581 ? 8'h10 : _T_4165; // @[Mux.scala 31:69:@2064.4]
  assign _T_4167 = _T_3578 ? 8'h8 : _T_4166; // @[Mux.scala 31:69:@2065.4]
  assign _T_4168 = _T_3575 ? 8'h4 : _T_4167; // @[Mux.scala 31:69:@2066.4]
  assign _T_4169 = _T_3572 ? 8'h2 : _T_4168; // @[Mux.scala 31:69:@2067.4]
  assign _T_4170 = _T_3569 ? 8'h1 : _T_4169; // @[Mux.scala 31:69:@2068.4]
  assign _T_4171 = _T_4170[0]; // @[OneHot.scala 66:30:@2069.4]
  assign _T_4172 = _T_4170[1]; // @[OneHot.scala 66:30:@2070.4]
  assign _T_4173 = _T_4170[2]; // @[OneHot.scala 66:30:@2071.4]
  assign _T_4174 = _T_4170[3]; // @[OneHot.scala 66:30:@2072.4]
  assign _T_4175 = _T_4170[4]; // @[OneHot.scala 66:30:@2073.4]
  assign _T_4176 = _T_4170[5]; // @[OneHot.scala 66:30:@2074.4]
  assign _T_4177 = _T_4170[6]; // @[OneHot.scala 66:30:@2075.4]
  assign _T_4178 = _T_4170[7]; // @[OneHot.scala 66:30:@2076.4]
  assign _T_4203 = _T_3569 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@2086.4]
  assign _T_4204 = _T_3590 ? 8'h40 : _T_4203; // @[Mux.scala 31:69:@2087.4]
  assign _T_4205 = _T_3587 ? 8'h20 : _T_4204; // @[Mux.scala 31:69:@2088.4]
  assign _T_4206 = _T_3584 ? 8'h10 : _T_4205; // @[Mux.scala 31:69:@2089.4]
  assign _T_4207 = _T_3581 ? 8'h8 : _T_4206; // @[Mux.scala 31:69:@2090.4]
  assign _T_4208 = _T_3578 ? 8'h4 : _T_4207; // @[Mux.scala 31:69:@2091.4]
  assign _T_4209 = _T_3575 ? 8'h2 : _T_4208; // @[Mux.scala 31:69:@2092.4]
  assign _T_4210 = _T_3572 ? 8'h1 : _T_4209; // @[Mux.scala 31:69:@2093.4]
  assign _T_4211 = _T_4210[0]; // @[OneHot.scala 66:30:@2094.4]
  assign _T_4212 = _T_4210[1]; // @[OneHot.scala 66:30:@2095.4]
  assign _T_4213 = _T_4210[2]; // @[OneHot.scala 66:30:@2096.4]
  assign _T_4214 = _T_4210[3]; // @[OneHot.scala 66:30:@2097.4]
  assign _T_4215 = _T_4210[4]; // @[OneHot.scala 66:30:@2098.4]
  assign _T_4216 = _T_4210[5]; // @[OneHot.scala 66:30:@2099.4]
  assign _T_4217 = _T_4210[6]; // @[OneHot.scala 66:30:@2100.4]
  assign _T_4218 = _T_4210[7]; // @[OneHot.scala 66:30:@2101.4]
  assign _T_4243 = _T_3572 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@2111.4]
  assign _T_4244 = _T_3569 ? 8'h40 : _T_4243; // @[Mux.scala 31:69:@2112.4]
  assign _T_4245 = _T_3590 ? 8'h20 : _T_4244; // @[Mux.scala 31:69:@2113.4]
  assign _T_4246 = _T_3587 ? 8'h10 : _T_4245; // @[Mux.scala 31:69:@2114.4]
  assign _T_4247 = _T_3584 ? 8'h8 : _T_4246; // @[Mux.scala 31:69:@2115.4]
  assign _T_4248 = _T_3581 ? 8'h4 : _T_4247; // @[Mux.scala 31:69:@2116.4]
  assign _T_4249 = _T_3578 ? 8'h2 : _T_4248; // @[Mux.scala 31:69:@2117.4]
  assign _T_4250 = _T_3575 ? 8'h1 : _T_4249; // @[Mux.scala 31:69:@2118.4]
  assign _T_4251 = _T_4250[0]; // @[OneHot.scala 66:30:@2119.4]
  assign _T_4252 = _T_4250[1]; // @[OneHot.scala 66:30:@2120.4]
  assign _T_4253 = _T_4250[2]; // @[OneHot.scala 66:30:@2121.4]
  assign _T_4254 = _T_4250[3]; // @[OneHot.scala 66:30:@2122.4]
  assign _T_4255 = _T_4250[4]; // @[OneHot.scala 66:30:@2123.4]
  assign _T_4256 = _T_4250[5]; // @[OneHot.scala 66:30:@2124.4]
  assign _T_4257 = _T_4250[6]; // @[OneHot.scala 66:30:@2125.4]
  assign _T_4258 = _T_4250[7]; // @[OneHot.scala 66:30:@2126.4]
  assign _T_4283 = _T_3575 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@2136.4]
  assign _T_4284 = _T_3572 ? 8'h40 : _T_4283; // @[Mux.scala 31:69:@2137.4]
  assign _T_4285 = _T_3569 ? 8'h20 : _T_4284; // @[Mux.scala 31:69:@2138.4]
  assign _T_4286 = _T_3590 ? 8'h10 : _T_4285; // @[Mux.scala 31:69:@2139.4]
  assign _T_4287 = _T_3587 ? 8'h8 : _T_4286; // @[Mux.scala 31:69:@2140.4]
  assign _T_4288 = _T_3584 ? 8'h4 : _T_4287; // @[Mux.scala 31:69:@2141.4]
  assign _T_4289 = _T_3581 ? 8'h2 : _T_4288; // @[Mux.scala 31:69:@2142.4]
  assign _T_4290 = _T_3578 ? 8'h1 : _T_4289; // @[Mux.scala 31:69:@2143.4]
  assign _T_4291 = _T_4290[0]; // @[OneHot.scala 66:30:@2144.4]
  assign _T_4292 = _T_4290[1]; // @[OneHot.scala 66:30:@2145.4]
  assign _T_4293 = _T_4290[2]; // @[OneHot.scala 66:30:@2146.4]
  assign _T_4294 = _T_4290[3]; // @[OneHot.scala 66:30:@2147.4]
  assign _T_4295 = _T_4290[4]; // @[OneHot.scala 66:30:@2148.4]
  assign _T_4296 = _T_4290[5]; // @[OneHot.scala 66:30:@2149.4]
  assign _T_4297 = _T_4290[6]; // @[OneHot.scala 66:30:@2150.4]
  assign _T_4298 = _T_4290[7]; // @[OneHot.scala 66:30:@2151.4]
  assign _T_4323 = _T_3578 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@2161.4]
  assign _T_4324 = _T_3575 ? 8'h40 : _T_4323; // @[Mux.scala 31:69:@2162.4]
  assign _T_4325 = _T_3572 ? 8'h20 : _T_4324; // @[Mux.scala 31:69:@2163.4]
  assign _T_4326 = _T_3569 ? 8'h10 : _T_4325; // @[Mux.scala 31:69:@2164.4]
  assign _T_4327 = _T_3590 ? 8'h8 : _T_4326; // @[Mux.scala 31:69:@2165.4]
  assign _T_4328 = _T_3587 ? 8'h4 : _T_4327; // @[Mux.scala 31:69:@2166.4]
  assign _T_4329 = _T_3584 ? 8'h2 : _T_4328; // @[Mux.scala 31:69:@2167.4]
  assign _T_4330 = _T_3581 ? 8'h1 : _T_4329; // @[Mux.scala 31:69:@2168.4]
  assign _T_4331 = _T_4330[0]; // @[OneHot.scala 66:30:@2169.4]
  assign _T_4332 = _T_4330[1]; // @[OneHot.scala 66:30:@2170.4]
  assign _T_4333 = _T_4330[2]; // @[OneHot.scala 66:30:@2171.4]
  assign _T_4334 = _T_4330[3]; // @[OneHot.scala 66:30:@2172.4]
  assign _T_4335 = _T_4330[4]; // @[OneHot.scala 66:30:@2173.4]
  assign _T_4336 = _T_4330[5]; // @[OneHot.scala 66:30:@2174.4]
  assign _T_4337 = _T_4330[6]; // @[OneHot.scala 66:30:@2175.4]
  assign _T_4338 = _T_4330[7]; // @[OneHot.scala 66:30:@2176.4]
  assign _T_4363 = _T_3581 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@2186.4]
  assign _T_4364 = _T_3578 ? 8'h40 : _T_4363; // @[Mux.scala 31:69:@2187.4]
  assign _T_4365 = _T_3575 ? 8'h20 : _T_4364; // @[Mux.scala 31:69:@2188.4]
  assign _T_4366 = _T_3572 ? 8'h10 : _T_4365; // @[Mux.scala 31:69:@2189.4]
  assign _T_4367 = _T_3569 ? 8'h8 : _T_4366; // @[Mux.scala 31:69:@2190.4]
  assign _T_4368 = _T_3590 ? 8'h4 : _T_4367; // @[Mux.scala 31:69:@2191.4]
  assign _T_4369 = _T_3587 ? 8'h2 : _T_4368; // @[Mux.scala 31:69:@2192.4]
  assign _T_4370 = _T_3584 ? 8'h1 : _T_4369; // @[Mux.scala 31:69:@2193.4]
  assign _T_4371 = _T_4370[0]; // @[OneHot.scala 66:30:@2194.4]
  assign _T_4372 = _T_4370[1]; // @[OneHot.scala 66:30:@2195.4]
  assign _T_4373 = _T_4370[2]; // @[OneHot.scala 66:30:@2196.4]
  assign _T_4374 = _T_4370[3]; // @[OneHot.scala 66:30:@2197.4]
  assign _T_4375 = _T_4370[4]; // @[OneHot.scala 66:30:@2198.4]
  assign _T_4376 = _T_4370[5]; // @[OneHot.scala 66:30:@2199.4]
  assign _T_4377 = _T_4370[6]; // @[OneHot.scala 66:30:@2200.4]
  assign _T_4378 = _T_4370[7]; // @[OneHot.scala 66:30:@2201.4]
  assign _T_4403 = _T_3584 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@2211.4]
  assign _T_4404 = _T_3581 ? 8'h40 : _T_4403; // @[Mux.scala 31:69:@2212.4]
  assign _T_4405 = _T_3578 ? 8'h20 : _T_4404; // @[Mux.scala 31:69:@2213.4]
  assign _T_4406 = _T_3575 ? 8'h10 : _T_4405; // @[Mux.scala 31:69:@2214.4]
  assign _T_4407 = _T_3572 ? 8'h8 : _T_4406; // @[Mux.scala 31:69:@2215.4]
  assign _T_4408 = _T_3569 ? 8'h4 : _T_4407; // @[Mux.scala 31:69:@2216.4]
  assign _T_4409 = _T_3590 ? 8'h2 : _T_4408; // @[Mux.scala 31:69:@2217.4]
  assign _T_4410 = _T_3587 ? 8'h1 : _T_4409; // @[Mux.scala 31:69:@2218.4]
  assign _T_4411 = _T_4410[0]; // @[OneHot.scala 66:30:@2219.4]
  assign _T_4412 = _T_4410[1]; // @[OneHot.scala 66:30:@2220.4]
  assign _T_4413 = _T_4410[2]; // @[OneHot.scala 66:30:@2221.4]
  assign _T_4414 = _T_4410[3]; // @[OneHot.scala 66:30:@2222.4]
  assign _T_4415 = _T_4410[4]; // @[OneHot.scala 66:30:@2223.4]
  assign _T_4416 = _T_4410[5]; // @[OneHot.scala 66:30:@2224.4]
  assign _T_4417 = _T_4410[6]; // @[OneHot.scala 66:30:@2225.4]
  assign _T_4418 = _T_4410[7]; // @[OneHot.scala 66:30:@2226.4]
  assign _T_4443 = _T_3587 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@2236.4]
  assign _T_4444 = _T_3584 ? 8'h40 : _T_4443; // @[Mux.scala 31:69:@2237.4]
  assign _T_4445 = _T_3581 ? 8'h20 : _T_4444; // @[Mux.scala 31:69:@2238.4]
  assign _T_4446 = _T_3578 ? 8'h10 : _T_4445; // @[Mux.scala 31:69:@2239.4]
  assign _T_4447 = _T_3575 ? 8'h8 : _T_4446; // @[Mux.scala 31:69:@2240.4]
  assign _T_4448 = _T_3572 ? 8'h4 : _T_4447; // @[Mux.scala 31:69:@2241.4]
  assign _T_4449 = _T_3569 ? 8'h2 : _T_4448; // @[Mux.scala 31:69:@2242.4]
  assign _T_4450 = _T_3590 ? 8'h1 : _T_4449; // @[Mux.scala 31:69:@2243.4]
  assign _T_4451 = _T_4450[0]; // @[OneHot.scala 66:30:@2244.4]
  assign _T_4452 = _T_4450[1]; // @[OneHot.scala 66:30:@2245.4]
  assign _T_4453 = _T_4450[2]; // @[OneHot.scala 66:30:@2246.4]
  assign _T_4454 = _T_4450[3]; // @[OneHot.scala 66:30:@2247.4]
  assign _T_4455 = _T_4450[4]; // @[OneHot.scala 66:30:@2248.4]
  assign _T_4456 = _T_4450[5]; // @[OneHot.scala 66:30:@2249.4]
  assign _T_4457 = _T_4450[6]; // @[OneHot.scala 66:30:@2250.4]
  assign _T_4458 = _T_4450[7]; // @[OneHot.scala 66:30:@2251.4]
  assign _T_4499 = {_T_4178,_T_4177,_T_4176,_T_4175,_T_4174,_T_4173,_T_4172,_T_4171}; // @[Mux.scala 19:72:@2267.4]
  assign _T_4501 = _T_2489 ? _T_4499 : 8'h0; // @[Mux.scala 19:72:@2268.4]
  assign _T_4508 = {_T_4217,_T_4216,_T_4215,_T_4214,_T_4213,_T_4212,_T_4211,_T_4218}; // @[Mux.scala 19:72:@2275.4]
  assign _T_4510 = _T_2490 ? _T_4508 : 8'h0; // @[Mux.scala 19:72:@2276.4]
  assign _T_4517 = {_T_4256,_T_4255,_T_4254,_T_4253,_T_4252,_T_4251,_T_4258,_T_4257}; // @[Mux.scala 19:72:@2283.4]
  assign _T_4519 = _T_2491 ? _T_4517 : 8'h0; // @[Mux.scala 19:72:@2284.4]
  assign _T_4526 = {_T_4295,_T_4294,_T_4293,_T_4292,_T_4291,_T_4298,_T_4297,_T_4296}; // @[Mux.scala 19:72:@2291.4]
  assign _T_4528 = _T_2492 ? _T_4526 : 8'h0; // @[Mux.scala 19:72:@2292.4]
  assign _T_4535 = {_T_4334,_T_4333,_T_4332,_T_4331,_T_4338,_T_4337,_T_4336,_T_4335}; // @[Mux.scala 19:72:@2299.4]
  assign _T_4537 = _T_2493 ? _T_4535 : 8'h0; // @[Mux.scala 19:72:@2300.4]
  assign _T_4544 = {_T_4373,_T_4372,_T_4371,_T_4378,_T_4377,_T_4376,_T_4375,_T_4374}; // @[Mux.scala 19:72:@2307.4]
  assign _T_4546 = _T_2494 ? _T_4544 : 8'h0; // @[Mux.scala 19:72:@2308.4]
  assign _T_4553 = {_T_4412,_T_4411,_T_4418,_T_4417,_T_4416,_T_4415,_T_4414,_T_4413}; // @[Mux.scala 19:72:@2315.4]
  assign _T_4555 = _T_2495 ? _T_4553 : 8'h0; // @[Mux.scala 19:72:@2316.4]
  assign _T_4562 = {_T_4451,_T_4458,_T_4457,_T_4456,_T_4455,_T_4454,_T_4453,_T_4452}; // @[Mux.scala 19:72:@2323.4]
  assign _T_4564 = _T_2496 ? _T_4562 : 8'h0; // @[Mux.scala 19:72:@2324.4]
  assign _T_4565 = _T_4501 | _T_4510; // @[Mux.scala 19:72:@2325.4]
  assign _T_4566 = _T_4565 | _T_4519; // @[Mux.scala 19:72:@2326.4]
  assign _T_4567 = _T_4566 | _T_4528; // @[Mux.scala 19:72:@2327.4]
  assign _T_4568 = _T_4567 | _T_4537; // @[Mux.scala 19:72:@2328.4]
  assign _T_4569 = _T_4568 | _T_4546; // @[Mux.scala 19:72:@2329.4]
  assign _T_4570 = _T_4569 | _T_4555; // @[Mux.scala 19:72:@2330.4]
  assign _T_4571 = _T_4570 | _T_4564; // @[Mux.scala 19:72:@2331.4]
  assign inputDataPriorityPorts_1_0 = _T_4571[0]; // @[Mux.scala 19:72:@2335.4]
  assign inputDataPriorityPorts_1_1 = _T_4571[1]; // @[Mux.scala 19:72:@2337.4]
  assign inputDataPriorityPorts_1_2 = _T_4571[2]; // @[Mux.scala 19:72:@2339.4]
  assign inputDataPriorityPorts_1_3 = _T_4571[3]; // @[Mux.scala 19:72:@2341.4]
  assign inputDataPriorityPorts_1_4 = _T_4571[4]; // @[Mux.scala 19:72:@2343.4]
  assign inputDataPriorityPorts_1_5 = _T_4571[5]; // @[Mux.scala 19:72:@2345.4]
  assign inputDataPriorityPorts_1_6 = _T_4571[6]; // @[Mux.scala 19:72:@2347.4]
  assign inputDataPriorityPorts_1_7 = _T_4571[7]; // @[Mux.scala 19:72:@2349.4]
  assign _T_4653 = inputAddrPriorityPorts_0_0 & _T_2410; // @[StoreQueue.scala 209:52:@2365.6]
  assign _T_4654 = _T_4653 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@2366.6]
  assign _T_4657 = inputAddrPriorityPorts_1_0 & _T_2410; // @[StoreQueue.scala 209:52:@2368.6]
  assign _T_4658 = _T_4657 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@2369.6]
  assign _T_4669 = _T_4654 | _T_4658; // @[StoreQueue.scala 210:30:@2374.6]
  assign _T_4670 = {_T_4658,_T_4654}; // @[OneHot.scala 18:45:@2376.8]
  assign _T_4671 = _T_4670[1]; // @[CircuitMath.scala 30:8:@2377.8]
  assign _GEN_305 = _T_4671 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@2378.8]
  assign _GEN_306 = _T_4669 ? _GEN_305 : addrQ_0; // @[StoreQueue.scala 210:40:@2375.6]
  assign _GEN_307 = _T_4669 ? 1'h1 : addrKnown_0; // @[StoreQueue.scala 210:40:@2375.6]
  assign _T_4676 = inputDataPriorityPorts_0_0 & _T_2448; // @[StoreQueue.scala 215:52:@2382.6]
  assign _T_4677 = _T_4676 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@2383.6]
  assign _T_4680 = inputDataPriorityPorts_1_0 & _T_2448; // @[StoreQueue.scala 215:52:@2385.6]
  assign _T_4681 = _T_4680 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@2386.6]
  assign _T_4692 = _T_4677 | _T_4681; // @[StoreQueue.scala 216:30:@2391.6]
  assign _T_4693 = {_T_4681,_T_4677}; // @[OneHot.scala 18:45:@2393.8]
  assign _T_4694 = _T_4693[1]; // @[CircuitMath.scala 30:8:@2394.8]
  assign _GEN_309 = _T_4694 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@2395.8]
  assign _GEN_310 = _T_4692 ? _GEN_309 : dataQ_0; // @[StoreQueue.scala 216:40:@2392.6]
  assign _GEN_311 = _T_4692 ? 1'h1 : dataKnown_0; // @[StoreQueue.scala 216:40:@2392.6]
  assign _GEN_312 = initBits_0 ? 1'h0 : _GEN_307; // @[StoreQueue.scala 204:35:@2359.4]
  assign _GEN_313 = initBits_0 ? 1'h0 : _GEN_311; // @[StoreQueue.scala 204:35:@2359.4]
  assign _GEN_314 = initBits_0 ? addrQ_0 : _GEN_306; // @[StoreQueue.scala 204:35:@2359.4]
  assign _GEN_315 = initBits_0 ? dataQ_0 : _GEN_310; // @[StoreQueue.scala 204:35:@2359.4]
  assign _T_4701 = inputAddrPriorityPorts_0_1 & _T_2413; // @[StoreQueue.scala 209:52:@2405.6]
  assign _T_4702 = _T_4701 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@2406.6]
  assign _T_4705 = inputAddrPriorityPorts_1_1 & _T_2413; // @[StoreQueue.scala 209:52:@2408.6]
  assign _T_4706 = _T_4705 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@2409.6]
  assign _T_4717 = _T_4702 | _T_4706; // @[StoreQueue.scala 210:30:@2414.6]
  assign _T_4718 = {_T_4706,_T_4702}; // @[OneHot.scala 18:45:@2416.8]
  assign _T_4719 = _T_4718[1]; // @[CircuitMath.scala 30:8:@2417.8]
  assign _GEN_317 = _T_4719 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@2418.8]
  assign _GEN_318 = _T_4717 ? _GEN_317 : addrQ_1; // @[StoreQueue.scala 210:40:@2415.6]
  assign _GEN_319 = _T_4717 ? 1'h1 : addrKnown_1; // @[StoreQueue.scala 210:40:@2415.6]
  assign _T_4724 = inputDataPriorityPorts_0_1 & _T_2451; // @[StoreQueue.scala 215:52:@2422.6]
  assign _T_4725 = _T_4724 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@2423.6]
  assign _T_4728 = inputDataPriorityPorts_1_1 & _T_2451; // @[StoreQueue.scala 215:52:@2425.6]
  assign _T_4729 = _T_4728 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@2426.6]
  assign _T_4740 = _T_4725 | _T_4729; // @[StoreQueue.scala 216:30:@2431.6]
  assign _T_4741 = {_T_4729,_T_4725}; // @[OneHot.scala 18:45:@2433.8]
  assign _T_4742 = _T_4741[1]; // @[CircuitMath.scala 30:8:@2434.8]
  assign _GEN_321 = _T_4742 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@2435.8]
  assign _GEN_322 = _T_4740 ? _GEN_321 : dataQ_1; // @[StoreQueue.scala 216:40:@2432.6]
  assign _GEN_323 = _T_4740 ? 1'h1 : dataKnown_1; // @[StoreQueue.scala 216:40:@2432.6]
  assign _GEN_324 = initBits_1 ? 1'h0 : _GEN_319; // @[StoreQueue.scala 204:35:@2399.4]
  assign _GEN_325 = initBits_1 ? 1'h0 : _GEN_323; // @[StoreQueue.scala 204:35:@2399.4]
  assign _GEN_326 = initBits_1 ? addrQ_1 : _GEN_318; // @[StoreQueue.scala 204:35:@2399.4]
  assign _GEN_327 = initBits_1 ? dataQ_1 : _GEN_322; // @[StoreQueue.scala 204:35:@2399.4]
  assign _T_4749 = inputAddrPriorityPorts_0_2 & _T_2416; // @[StoreQueue.scala 209:52:@2445.6]
  assign _T_4750 = _T_4749 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@2446.6]
  assign _T_4753 = inputAddrPriorityPorts_1_2 & _T_2416; // @[StoreQueue.scala 209:52:@2448.6]
  assign _T_4754 = _T_4753 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@2449.6]
  assign _T_4765 = _T_4750 | _T_4754; // @[StoreQueue.scala 210:30:@2454.6]
  assign _T_4766 = {_T_4754,_T_4750}; // @[OneHot.scala 18:45:@2456.8]
  assign _T_4767 = _T_4766[1]; // @[CircuitMath.scala 30:8:@2457.8]
  assign _GEN_329 = _T_4767 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@2458.8]
  assign _GEN_330 = _T_4765 ? _GEN_329 : addrQ_2; // @[StoreQueue.scala 210:40:@2455.6]
  assign _GEN_331 = _T_4765 ? 1'h1 : addrKnown_2; // @[StoreQueue.scala 210:40:@2455.6]
  assign _T_4772 = inputDataPriorityPorts_0_2 & _T_2454; // @[StoreQueue.scala 215:52:@2462.6]
  assign _T_4773 = _T_4772 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@2463.6]
  assign _T_4776 = inputDataPriorityPorts_1_2 & _T_2454; // @[StoreQueue.scala 215:52:@2465.6]
  assign _T_4777 = _T_4776 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@2466.6]
  assign _T_4788 = _T_4773 | _T_4777; // @[StoreQueue.scala 216:30:@2471.6]
  assign _T_4789 = {_T_4777,_T_4773}; // @[OneHot.scala 18:45:@2473.8]
  assign _T_4790 = _T_4789[1]; // @[CircuitMath.scala 30:8:@2474.8]
  assign _GEN_333 = _T_4790 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@2475.8]
  assign _GEN_334 = _T_4788 ? _GEN_333 : dataQ_2; // @[StoreQueue.scala 216:40:@2472.6]
  assign _GEN_335 = _T_4788 ? 1'h1 : dataKnown_2; // @[StoreQueue.scala 216:40:@2472.6]
  assign _GEN_336 = initBits_2 ? 1'h0 : _GEN_331; // @[StoreQueue.scala 204:35:@2439.4]
  assign _GEN_337 = initBits_2 ? 1'h0 : _GEN_335; // @[StoreQueue.scala 204:35:@2439.4]
  assign _GEN_338 = initBits_2 ? addrQ_2 : _GEN_330; // @[StoreQueue.scala 204:35:@2439.4]
  assign _GEN_339 = initBits_2 ? dataQ_2 : _GEN_334; // @[StoreQueue.scala 204:35:@2439.4]
  assign _T_4797 = inputAddrPriorityPorts_0_3 & _T_2419; // @[StoreQueue.scala 209:52:@2485.6]
  assign _T_4798 = _T_4797 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@2486.6]
  assign _T_4801 = inputAddrPriorityPorts_1_3 & _T_2419; // @[StoreQueue.scala 209:52:@2488.6]
  assign _T_4802 = _T_4801 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@2489.6]
  assign _T_4813 = _T_4798 | _T_4802; // @[StoreQueue.scala 210:30:@2494.6]
  assign _T_4814 = {_T_4802,_T_4798}; // @[OneHot.scala 18:45:@2496.8]
  assign _T_4815 = _T_4814[1]; // @[CircuitMath.scala 30:8:@2497.8]
  assign _GEN_341 = _T_4815 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@2498.8]
  assign _GEN_342 = _T_4813 ? _GEN_341 : addrQ_3; // @[StoreQueue.scala 210:40:@2495.6]
  assign _GEN_343 = _T_4813 ? 1'h1 : addrKnown_3; // @[StoreQueue.scala 210:40:@2495.6]
  assign _T_4820 = inputDataPriorityPorts_0_3 & _T_2457; // @[StoreQueue.scala 215:52:@2502.6]
  assign _T_4821 = _T_4820 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@2503.6]
  assign _T_4824 = inputDataPriorityPorts_1_3 & _T_2457; // @[StoreQueue.scala 215:52:@2505.6]
  assign _T_4825 = _T_4824 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@2506.6]
  assign _T_4836 = _T_4821 | _T_4825; // @[StoreQueue.scala 216:30:@2511.6]
  assign _T_4837 = {_T_4825,_T_4821}; // @[OneHot.scala 18:45:@2513.8]
  assign _T_4838 = _T_4837[1]; // @[CircuitMath.scala 30:8:@2514.8]
  assign _GEN_345 = _T_4838 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@2515.8]
  assign _GEN_346 = _T_4836 ? _GEN_345 : dataQ_3; // @[StoreQueue.scala 216:40:@2512.6]
  assign _GEN_347 = _T_4836 ? 1'h1 : dataKnown_3; // @[StoreQueue.scala 216:40:@2512.6]
  assign _GEN_348 = initBits_3 ? 1'h0 : _GEN_343; // @[StoreQueue.scala 204:35:@2479.4]
  assign _GEN_349 = initBits_3 ? 1'h0 : _GEN_347; // @[StoreQueue.scala 204:35:@2479.4]
  assign _GEN_350 = initBits_3 ? addrQ_3 : _GEN_342; // @[StoreQueue.scala 204:35:@2479.4]
  assign _GEN_351 = initBits_3 ? dataQ_3 : _GEN_346; // @[StoreQueue.scala 204:35:@2479.4]
  assign _T_4845 = inputAddrPriorityPorts_0_4 & _T_2422; // @[StoreQueue.scala 209:52:@2525.6]
  assign _T_4846 = _T_4845 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@2526.6]
  assign _T_4849 = inputAddrPriorityPorts_1_4 & _T_2422; // @[StoreQueue.scala 209:52:@2528.6]
  assign _T_4850 = _T_4849 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@2529.6]
  assign _T_4861 = _T_4846 | _T_4850; // @[StoreQueue.scala 210:30:@2534.6]
  assign _T_4862 = {_T_4850,_T_4846}; // @[OneHot.scala 18:45:@2536.8]
  assign _T_4863 = _T_4862[1]; // @[CircuitMath.scala 30:8:@2537.8]
  assign _GEN_353 = _T_4863 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@2538.8]
  assign _GEN_354 = _T_4861 ? _GEN_353 : addrQ_4; // @[StoreQueue.scala 210:40:@2535.6]
  assign _GEN_355 = _T_4861 ? 1'h1 : addrKnown_4; // @[StoreQueue.scala 210:40:@2535.6]
  assign _T_4868 = inputDataPriorityPorts_0_4 & _T_2460; // @[StoreQueue.scala 215:52:@2542.6]
  assign _T_4869 = _T_4868 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@2543.6]
  assign _T_4872 = inputDataPriorityPorts_1_4 & _T_2460; // @[StoreQueue.scala 215:52:@2545.6]
  assign _T_4873 = _T_4872 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@2546.6]
  assign _T_4884 = _T_4869 | _T_4873; // @[StoreQueue.scala 216:30:@2551.6]
  assign _T_4885 = {_T_4873,_T_4869}; // @[OneHot.scala 18:45:@2553.8]
  assign _T_4886 = _T_4885[1]; // @[CircuitMath.scala 30:8:@2554.8]
  assign _GEN_357 = _T_4886 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@2555.8]
  assign _GEN_358 = _T_4884 ? _GEN_357 : dataQ_4; // @[StoreQueue.scala 216:40:@2552.6]
  assign _GEN_359 = _T_4884 ? 1'h1 : dataKnown_4; // @[StoreQueue.scala 216:40:@2552.6]
  assign _GEN_360 = initBits_4 ? 1'h0 : _GEN_355; // @[StoreQueue.scala 204:35:@2519.4]
  assign _GEN_361 = initBits_4 ? 1'h0 : _GEN_359; // @[StoreQueue.scala 204:35:@2519.4]
  assign _GEN_362 = initBits_4 ? addrQ_4 : _GEN_354; // @[StoreQueue.scala 204:35:@2519.4]
  assign _GEN_363 = initBits_4 ? dataQ_4 : _GEN_358; // @[StoreQueue.scala 204:35:@2519.4]
  assign _T_4893 = inputAddrPriorityPorts_0_5 & _T_2425; // @[StoreQueue.scala 209:52:@2565.6]
  assign _T_4894 = _T_4893 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@2566.6]
  assign _T_4897 = inputAddrPriorityPorts_1_5 & _T_2425; // @[StoreQueue.scala 209:52:@2568.6]
  assign _T_4898 = _T_4897 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@2569.6]
  assign _T_4909 = _T_4894 | _T_4898; // @[StoreQueue.scala 210:30:@2574.6]
  assign _T_4910 = {_T_4898,_T_4894}; // @[OneHot.scala 18:45:@2576.8]
  assign _T_4911 = _T_4910[1]; // @[CircuitMath.scala 30:8:@2577.8]
  assign _GEN_365 = _T_4911 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@2578.8]
  assign _GEN_366 = _T_4909 ? _GEN_365 : addrQ_5; // @[StoreQueue.scala 210:40:@2575.6]
  assign _GEN_367 = _T_4909 ? 1'h1 : addrKnown_5; // @[StoreQueue.scala 210:40:@2575.6]
  assign _T_4916 = inputDataPriorityPorts_0_5 & _T_2463; // @[StoreQueue.scala 215:52:@2582.6]
  assign _T_4917 = _T_4916 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@2583.6]
  assign _T_4920 = inputDataPriorityPorts_1_5 & _T_2463; // @[StoreQueue.scala 215:52:@2585.6]
  assign _T_4921 = _T_4920 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@2586.6]
  assign _T_4932 = _T_4917 | _T_4921; // @[StoreQueue.scala 216:30:@2591.6]
  assign _T_4933 = {_T_4921,_T_4917}; // @[OneHot.scala 18:45:@2593.8]
  assign _T_4934 = _T_4933[1]; // @[CircuitMath.scala 30:8:@2594.8]
  assign _GEN_369 = _T_4934 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@2595.8]
  assign _GEN_370 = _T_4932 ? _GEN_369 : dataQ_5; // @[StoreQueue.scala 216:40:@2592.6]
  assign _GEN_371 = _T_4932 ? 1'h1 : dataKnown_5; // @[StoreQueue.scala 216:40:@2592.6]
  assign _GEN_372 = initBits_5 ? 1'h0 : _GEN_367; // @[StoreQueue.scala 204:35:@2559.4]
  assign _GEN_373 = initBits_5 ? 1'h0 : _GEN_371; // @[StoreQueue.scala 204:35:@2559.4]
  assign _GEN_374 = initBits_5 ? addrQ_5 : _GEN_366; // @[StoreQueue.scala 204:35:@2559.4]
  assign _GEN_375 = initBits_5 ? dataQ_5 : _GEN_370; // @[StoreQueue.scala 204:35:@2559.4]
  assign _T_4941 = inputAddrPriorityPorts_0_6 & _T_2428; // @[StoreQueue.scala 209:52:@2605.6]
  assign _T_4942 = _T_4941 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@2606.6]
  assign _T_4945 = inputAddrPriorityPorts_1_6 & _T_2428; // @[StoreQueue.scala 209:52:@2608.6]
  assign _T_4946 = _T_4945 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@2609.6]
  assign _T_4957 = _T_4942 | _T_4946; // @[StoreQueue.scala 210:30:@2614.6]
  assign _T_4958 = {_T_4946,_T_4942}; // @[OneHot.scala 18:45:@2616.8]
  assign _T_4959 = _T_4958[1]; // @[CircuitMath.scala 30:8:@2617.8]
  assign _GEN_377 = _T_4959 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@2618.8]
  assign _GEN_378 = _T_4957 ? _GEN_377 : addrQ_6; // @[StoreQueue.scala 210:40:@2615.6]
  assign _GEN_379 = _T_4957 ? 1'h1 : addrKnown_6; // @[StoreQueue.scala 210:40:@2615.6]
  assign _T_4964 = inputDataPriorityPorts_0_6 & _T_2466; // @[StoreQueue.scala 215:52:@2622.6]
  assign _T_4965 = _T_4964 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@2623.6]
  assign _T_4968 = inputDataPriorityPorts_1_6 & _T_2466; // @[StoreQueue.scala 215:52:@2625.6]
  assign _T_4969 = _T_4968 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@2626.6]
  assign _T_4980 = _T_4965 | _T_4969; // @[StoreQueue.scala 216:30:@2631.6]
  assign _T_4981 = {_T_4969,_T_4965}; // @[OneHot.scala 18:45:@2633.8]
  assign _T_4982 = _T_4981[1]; // @[CircuitMath.scala 30:8:@2634.8]
  assign _GEN_381 = _T_4982 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@2635.8]
  assign _GEN_382 = _T_4980 ? _GEN_381 : dataQ_6; // @[StoreQueue.scala 216:40:@2632.6]
  assign _GEN_383 = _T_4980 ? 1'h1 : dataKnown_6; // @[StoreQueue.scala 216:40:@2632.6]
  assign _GEN_384 = initBits_6 ? 1'h0 : _GEN_379; // @[StoreQueue.scala 204:35:@2599.4]
  assign _GEN_385 = initBits_6 ? 1'h0 : _GEN_383; // @[StoreQueue.scala 204:35:@2599.4]
  assign _GEN_386 = initBits_6 ? addrQ_6 : _GEN_378; // @[StoreQueue.scala 204:35:@2599.4]
  assign _GEN_387 = initBits_6 ? dataQ_6 : _GEN_382; // @[StoreQueue.scala 204:35:@2599.4]
  assign _T_4989 = inputAddrPriorityPorts_0_7 & _T_2431; // @[StoreQueue.scala 209:52:@2645.6]
  assign _T_4990 = _T_4989 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@2646.6]
  assign _T_4993 = inputAddrPriorityPorts_1_7 & _T_2431; // @[StoreQueue.scala 209:52:@2648.6]
  assign _T_4994 = _T_4993 & io_storeAddrEnable_1; // @[StoreQueue.scala 209:81:@2649.6]
  assign _T_5005 = _T_4990 | _T_4994; // @[StoreQueue.scala 210:30:@2654.6]
  assign _T_5006 = {_T_4994,_T_4990}; // @[OneHot.scala 18:45:@2656.8]
  assign _T_5007 = _T_5006[1]; // @[CircuitMath.scala 30:8:@2657.8]
  assign _GEN_389 = _T_5007 ? io_addressFromStorePorts_1 : io_addressFromStorePorts_0; // @[StoreQueue.scala 211:30:@2658.8]
  assign _GEN_390 = _T_5005 ? _GEN_389 : addrQ_7; // @[StoreQueue.scala 210:40:@2655.6]
  assign _GEN_391 = _T_5005 ? 1'h1 : addrKnown_7; // @[StoreQueue.scala 210:40:@2655.6]
  assign _T_5012 = inputDataPriorityPorts_0_7 & _T_2469; // @[StoreQueue.scala 215:52:@2662.6]
  assign _T_5013 = _T_5012 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@2663.6]
  assign _T_5016 = inputDataPriorityPorts_1_7 & _T_2469; // @[StoreQueue.scala 215:52:@2665.6]
  assign _T_5017 = _T_5016 & io_storeDataEnable_1; // @[StoreQueue.scala 215:81:@2666.6]
  assign _T_5028 = _T_5013 | _T_5017; // @[StoreQueue.scala 216:30:@2671.6]
  assign _T_5029 = {_T_5017,_T_5013}; // @[OneHot.scala 18:45:@2673.8]
  assign _T_5030 = _T_5029[1]; // @[CircuitMath.scala 30:8:@2674.8]
  assign _GEN_393 = _T_5030 ? io_dataFromStorePorts_1 : io_dataFromStorePorts_0; // @[StoreQueue.scala 217:30:@2675.8]
  assign _GEN_394 = _T_5028 ? _GEN_393 : dataQ_7; // @[StoreQueue.scala 216:40:@2672.6]
  assign _GEN_395 = _T_5028 ? 1'h1 : dataKnown_7; // @[StoreQueue.scala 216:40:@2672.6]
  assign _GEN_396 = initBits_7 ? 1'h0 : _GEN_391; // @[StoreQueue.scala 204:35:@2639.4]
  assign _GEN_397 = initBits_7 ? 1'h0 : _GEN_395; // @[StoreQueue.scala 204:35:@2639.4]
  assign _GEN_398 = initBits_7 ? addrQ_7 : _GEN_390; // @[StoreQueue.scala 204:35:@2639.4]
  assign _GEN_399 = initBits_7 ? dataQ_7 : _GEN_394; // @[StoreQueue.scala 204:35:@2639.4]
  assign _T_5033 = storeRequest & io_memIsReadyForStores; // @[StoreQueue.scala 229:23:@2679.4]
  assign _T_5036 = head + 3'h1; // @[util.scala 10:8:@2681.6]
  assign _GEN_144 = _T_5036 % 4'h8; // @[util.scala 10:14:@2682.6]
  assign _T_5037 = _GEN_144[3:0]; // @[util.scala 10:14:@2682.6]
  assign _GEN_400 = _T_5033 ? _T_5037 : {{1'd0}, head}; // @[StoreQueue.scala 229:50:@2680.4]
  assign _GEN_458 = {{1'd0}, io_bbNumStores}; // @[util.scala 10:8:@2686.6]
  assign _T_5039 = tail + _GEN_458; // @[util.scala 10:8:@2686.6]
  assign _GEN_145 = _T_5039 % 4'h8; // @[util.scala 10:14:@2687.6]
  assign _T_5040 = _GEN_145[3:0]; // @[util.scala 10:14:@2687.6]
  assign _GEN_401 = io_bbStart ? _T_5040 : {{1'd0}, tail}; // @[StoreQueue.scala 233:20:@2685.4]
  assign _T_5042 = allocatedEntries_0 == 1'h0; // @[StoreQueue.scala 237:84:@2690.4]
  assign _T_5043 = storeCompleted_0 | _T_5042; // @[StoreQueue.scala 237:81:@2691.4]
  assign _T_5045 = allocatedEntries_1 == 1'h0; // @[StoreQueue.scala 237:84:@2692.4]
  assign _T_5046 = storeCompleted_1 | _T_5045; // @[StoreQueue.scala 237:81:@2693.4]
  assign _T_5048 = allocatedEntries_2 == 1'h0; // @[StoreQueue.scala 237:84:@2694.4]
  assign _T_5049 = storeCompleted_2 | _T_5048; // @[StoreQueue.scala 237:81:@2695.4]
  assign _T_5051 = allocatedEntries_3 == 1'h0; // @[StoreQueue.scala 237:84:@2696.4]
  assign _T_5052 = storeCompleted_3 | _T_5051; // @[StoreQueue.scala 237:81:@2697.4]
  assign _T_5054 = allocatedEntries_4 == 1'h0; // @[StoreQueue.scala 237:84:@2698.4]
  assign _T_5055 = storeCompleted_4 | _T_5054; // @[StoreQueue.scala 237:81:@2699.4]
  assign _T_5057 = allocatedEntries_5 == 1'h0; // @[StoreQueue.scala 237:84:@2700.4]
  assign _T_5058 = storeCompleted_5 | _T_5057; // @[StoreQueue.scala 237:81:@2701.4]
  assign _T_5060 = allocatedEntries_6 == 1'h0; // @[StoreQueue.scala 237:84:@2702.4]
  assign _T_5061 = storeCompleted_6 | _T_5060; // @[StoreQueue.scala 237:81:@2703.4]
  assign _T_5063 = allocatedEntries_7 == 1'h0; // @[StoreQueue.scala 237:84:@2704.4]
  assign _T_5064 = storeCompleted_7 | _T_5063; // @[StoreQueue.scala 237:81:@2705.4]
  assign _T_5081 = _T_5043 & _T_5046; // @[StoreQueue.scala 237:98:@2716.4]
  assign _T_5082 = _T_5081 & _T_5049; // @[StoreQueue.scala 237:98:@2717.4]
  assign _T_5083 = _T_5082 & _T_5052; // @[StoreQueue.scala 237:98:@2718.4]
  assign _T_5084 = _T_5083 & _T_5055; // @[StoreQueue.scala 237:98:@2719.4]
  assign _T_5085 = _T_5084 & _T_5058; // @[StoreQueue.scala 237:98:@2720.4]
  assign _T_5086 = _T_5085 & _T_5061; // @[StoreQueue.scala 237:98:@2721.4]
  assign _GEN_403 = 3'h1 == head ? dataQ_1 : dataQ_0; // @[StoreQueue.scala 252:21:@2759.4]
  assign _GEN_404 = 3'h2 == head ? dataQ_2 : _GEN_403; // @[StoreQueue.scala 252:21:@2759.4]
  assign _GEN_405 = 3'h3 == head ? dataQ_3 : _GEN_404; // @[StoreQueue.scala 252:21:@2759.4]
  assign _GEN_406 = 3'h4 == head ? dataQ_4 : _GEN_405; // @[StoreQueue.scala 252:21:@2759.4]
  assign _GEN_407 = 3'h5 == head ? dataQ_5 : _GEN_406; // @[StoreQueue.scala 252:21:@2759.4]
  assign _GEN_408 = 3'h6 == head ? dataQ_6 : _GEN_407; // @[StoreQueue.scala 252:21:@2759.4]
  assign io_storeTail = tail; // @[StoreQueue.scala 246:16:@2725.4]
  assign io_storeHead = head; // @[StoreQueue.scala 245:16:@2724.4]
  assign io_storeEmpty = _T_5086 & _T_5064; // @[StoreQueue.scala 237:17:@2723.4]
  assign io_storeAddrDone_0 = addrKnown_0; // @[StoreQueue.scala 250:20:@2750.4]
  assign io_storeAddrDone_1 = addrKnown_1; // @[StoreQueue.scala 250:20:@2751.4]
  assign io_storeAddrDone_2 = addrKnown_2; // @[StoreQueue.scala 250:20:@2752.4]
  assign io_storeAddrDone_3 = addrKnown_3; // @[StoreQueue.scala 250:20:@2753.4]
  assign io_storeAddrDone_4 = addrKnown_4; // @[StoreQueue.scala 250:20:@2754.4]
  assign io_storeAddrDone_5 = addrKnown_5; // @[StoreQueue.scala 250:20:@2755.4]
  assign io_storeAddrDone_6 = addrKnown_6; // @[StoreQueue.scala 250:20:@2756.4]
  assign io_storeAddrDone_7 = addrKnown_7; // @[StoreQueue.scala 250:20:@2757.4]
  assign io_storeDataDone_0 = dataKnown_0; // @[StoreQueue.scala 249:20:@2742.4]
  assign io_storeDataDone_1 = dataKnown_1; // @[StoreQueue.scala 249:20:@2743.4]
  assign io_storeDataDone_2 = dataKnown_2; // @[StoreQueue.scala 249:20:@2744.4]
  assign io_storeDataDone_3 = dataKnown_3; // @[StoreQueue.scala 249:20:@2745.4]
  assign io_storeDataDone_4 = dataKnown_4; // @[StoreQueue.scala 249:20:@2746.4]
  assign io_storeDataDone_5 = dataKnown_5; // @[StoreQueue.scala 249:20:@2747.4]
  assign io_storeDataDone_6 = dataKnown_6; // @[StoreQueue.scala 249:20:@2748.4]
  assign io_storeDataDone_7 = dataKnown_7; // @[StoreQueue.scala 249:20:@2749.4]
  assign io_storeAddrQueue_0 = addrQ_0; // @[StoreQueue.scala 247:21:@2726.4]
  assign io_storeAddrQueue_1 = addrQ_1; // @[StoreQueue.scala 247:21:@2727.4]
  assign io_storeAddrQueue_2 = addrQ_2; // @[StoreQueue.scala 247:21:@2728.4]
  assign io_storeAddrQueue_3 = addrQ_3; // @[StoreQueue.scala 247:21:@2729.4]
  assign io_storeAddrQueue_4 = addrQ_4; // @[StoreQueue.scala 247:21:@2730.4]
  assign io_storeAddrQueue_5 = addrQ_5; // @[StoreQueue.scala 247:21:@2731.4]
  assign io_storeAddrQueue_6 = addrQ_6; // @[StoreQueue.scala 247:21:@2732.4]
  assign io_storeAddrQueue_7 = addrQ_7; // @[StoreQueue.scala 247:21:@2733.4]
  assign io_storeDataQueue_0 = dataQ_0; // @[StoreQueue.scala 248:21:@2734.4]
  assign io_storeDataQueue_1 = dataQ_1; // @[StoreQueue.scala 248:21:@2735.4]
  assign io_storeDataQueue_2 = dataQ_2; // @[StoreQueue.scala 248:21:@2736.4]
  assign io_storeDataQueue_3 = dataQ_3; // @[StoreQueue.scala 248:21:@2737.4]
  assign io_storeDataQueue_4 = dataQ_4; // @[StoreQueue.scala 248:21:@2738.4]
  assign io_storeDataQueue_5 = dataQ_5; // @[StoreQueue.scala 248:21:@2739.4]
  assign io_storeDataQueue_6 = dataQ_6; // @[StoreQueue.scala 248:21:@2740.4]
  assign io_storeDataQueue_7 = dataQ_7; // @[StoreQueue.scala 248:21:@2741.4]
  assign io_storeAddrToMem = 3'h7 == head ? addrQ_7 : _GEN_262; // @[StoreQueue.scala 253:21:@2760.4]
  assign io_storeDataToMem = 3'h7 == head ? dataQ_7 : _GEN_408; // @[StoreQueue.scala 252:21:@2759.4]
  assign io_storeEnableToMem = _T_1941 & _T_1950; // @[StoreQueue.scala 251:23:@2758.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  portQ_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  portQ_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  portQ_2 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  portQ_3 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  portQ_4 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  portQ_5 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  portQ_6 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  portQ_7 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  addrQ_0 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  addrQ_1 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  addrQ_2 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  addrQ_3 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  addrQ_4 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  addrQ_5 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  addrQ_6 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  addrQ_7 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  dataQ_0 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  dataQ_1 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  dataQ_2 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  dataQ_3 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  dataQ_4 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  dataQ_5 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  dataQ_6 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  dataQ_7 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrKnown_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrKnown_1 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrKnown_2 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrKnown_3 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrKnown_4 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrKnown_5 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrKnown_6 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrKnown_7 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  dataKnown_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  dataKnown_1 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  dataKnown_2 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  dataKnown_3 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  dataKnown_4 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  dataKnown_5 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  dataKnown_6 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  dataKnown_7 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  storeCompleted_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  storeCompleted_1 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  storeCompleted_2 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  storeCompleted_3 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  storeCompleted_4 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  storeCompleted_5 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  storeCompleted_6 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  storeCompleted_7 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  checkBits_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  checkBits_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  checkBits_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  checkBits_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  checkBits_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  checkBits_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  checkBits_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  checkBits_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  previousLoadHead = _RAND_74[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 3'h0;
    end else begin
      head <= _GEN_400[2:0];
    end
    if (reset) begin
      tail <= 3'h0;
    end else begin
      tail <= _GEN_401[2:0];
    end
    if (reset) begin
      offsetQ_0 <= 3'h0;
    end else begin
      if (initBits_0) begin
        if (3'h7 == _T_1068) begin
          offsetQ_0 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1068) begin
            offsetQ_0 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1068) begin
              offsetQ_0 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1068) begin
                offsetQ_0 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1068) begin
                  offsetQ_0 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1068) begin
                    offsetQ_0 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1068) begin
                      offsetQ_0 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_0 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 3'h0;
    end else begin
      if (initBits_1) begin
        if (3'h7 == _T_1086) begin
          offsetQ_1 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1086) begin
            offsetQ_1 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1086) begin
              offsetQ_1 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1086) begin
                offsetQ_1 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1086) begin
                  offsetQ_1 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1086) begin
                    offsetQ_1 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1086) begin
                      offsetQ_1 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_1 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 3'h0;
    end else begin
      if (initBits_2) begin
        if (3'h7 == _T_1104) begin
          offsetQ_2 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1104) begin
            offsetQ_2 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1104) begin
              offsetQ_2 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1104) begin
                offsetQ_2 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1104) begin
                  offsetQ_2 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1104) begin
                    offsetQ_2 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1104) begin
                      offsetQ_2 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_2 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 3'h0;
    end else begin
      if (initBits_3) begin
        if (3'h7 == _T_1122) begin
          offsetQ_3 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1122) begin
            offsetQ_3 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1122) begin
              offsetQ_3 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1122) begin
                offsetQ_3 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1122) begin
                  offsetQ_3 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1122) begin
                    offsetQ_3 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1122) begin
                      offsetQ_3 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_3 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 3'h0;
    end else begin
      if (initBits_4) begin
        if (3'h7 == _T_1140) begin
          offsetQ_4 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1140) begin
            offsetQ_4 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1140) begin
              offsetQ_4 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1140) begin
                offsetQ_4 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1140) begin
                  offsetQ_4 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1140) begin
                    offsetQ_4 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1140) begin
                      offsetQ_4 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_4 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 3'h0;
    end else begin
      if (initBits_5) begin
        if (3'h7 == _T_1158) begin
          offsetQ_5 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1158) begin
            offsetQ_5 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1158) begin
              offsetQ_5 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1158) begin
                offsetQ_5 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1158) begin
                  offsetQ_5 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1158) begin
                    offsetQ_5 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1158) begin
                      offsetQ_5 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_5 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 3'h0;
    end else begin
      if (initBits_6) begin
        if (3'h7 == _T_1176) begin
          offsetQ_6 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1176) begin
            offsetQ_6 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1176) begin
              offsetQ_6 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1176) begin
                offsetQ_6 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1176) begin
                  offsetQ_6 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1176) begin
                    offsetQ_6 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1176) begin
                      offsetQ_6 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_6 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 3'h0;
    end else begin
      if (initBits_7) begin
        if (3'h7 == _T_1194) begin
          offsetQ_7 <= io_bbStoreOffsets_7;
        end else begin
          if (3'h6 == _T_1194) begin
            offsetQ_7 <= io_bbStoreOffsets_6;
          end else begin
            if (3'h5 == _T_1194) begin
              offsetQ_7 <= io_bbStoreOffsets_5;
            end else begin
              if (3'h4 == _T_1194) begin
                offsetQ_7 <= io_bbStoreOffsets_4;
              end else begin
                if (3'h3 == _T_1194) begin
                  offsetQ_7 <= io_bbStoreOffsets_3;
                end else begin
                  if (3'h2 == _T_1194) begin
                    offsetQ_7 <= io_bbStoreOffsets_2;
                  end else begin
                    if (3'h1 == _T_1194) begin
                      offsetQ_7 <= io_bbStoreOffsets_1;
                    end else begin
                      offsetQ_7 <= io_bbStoreOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        if (3'h7 == _T_1068) begin
          portQ_0 <= 1'h0;
        end else begin
          if (3'h6 == _T_1068) begin
            portQ_0 <= 1'h0;
          end else begin
            if (3'h5 == _T_1068) begin
              portQ_0 <= 1'h0;
            end else begin
              if (3'h4 == _T_1068) begin
                portQ_0 <= 1'h0;
              end else begin
                if (3'h3 == _T_1068) begin
                  portQ_0 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1068) begin
                    portQ_0 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1068) begin
                      portQ_0 <= io_bbStorePorts_1;
                    end else begin
                      portQ_0 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        if (3'h7 == _T_1086) begin
          portQ_1 <= 1'h0;
        end else begin
          if (3'h6 == _T_1086) begin
            portQ_1 <= 1'h0;
          end else begin
            if (3'h5 == _T_1086) begin
              portQ_1 <= 1'h0;
            end else begin
              if (3'h4 == _T_1086) begin
                portQ_1 <= 1'h0;
              end else begin
                if (3'h3 == _T_1086) begin
                  portQ_1 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1086) begin
                    portQ_1 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1086) begin
                      portQ_1 <= io_bbStorePorts_1;
                    end else begin
                      portQ_1 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        if (3'h7 == _T_1104) begin
          portQ_2 <= 1'h0;
        end else begin
          if (3'h6 == _T_1104) begin
            portQ_2 <= 1'h0;
          end else begin
            if (3'h5 == _T_1104) begin
              portQ_2 <= 1'h0;
            end else begin
              if (3'h4 == _T_1104) begin
                portQ_2 <= 1'h0;
              end else begin
                if (3'h3 == _T_1104) begin
                  portQ_2 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1104) begin
                    portQ_2 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1104) begin
                      portQ_2 <= io_bbStorePorts_1;
                    end else begin
                      portQ_2 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        if (3'h7 == _T_1122) begin
          portQ_3 <= 1'h0;
        end else begin
          if (3'h6 == _T_1122) begin
            portQ_3 <= 1'h0;
          end else begin
            if (3'h5 == _T_1122) begin
              portQ_3 <= 1'h0;
            end else begin
              if (3'h4 == _T_1122) begin
                portQ_3 <= 1'h0;
              end else begin
                if (3'h3 == _T_1122) begin
                  portQ_3 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1122) begin
                    portQ_3 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1122) begin
                      portQ_3 <= io_bbStorePorts_1;
                    end else begin
                      portQ_3 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        if (3'h7 == _T_1140) begin
          portQ_4 <= 1'h0;
        end else begin
          if (3'h6 == _T_1140) begin
            portQ_4 <= 1'h0;
          end else begin
            if (3'h5 == _T_1140) begin
              portQ_4 <= 1'h0;
            end else begin
              if (3'h4 == _T_1140) begin
                portQ_4 <= 1'h0;
              end else begin
                if (3'h3 == _T_1140) begin
                  portQ_4 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1140) begin
                    portQ_4 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1140) begin
                      portQ_4 <= io_bbStorePorts_1;
                    end else begin
                      portQ_4 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        if (3'h7 == _T_1158) begin
          portQ_5 <= 1'h0;
        end else begin
          if (3'h6 == _T_1158) begin
            portQ_5 <= 1'h0;
          end else begin
            if (3'h5 == _T_1158) begin
              portQ_5 <= 1'h0;
            end else begin
              if (3'h4 == _T_1158) begin
                portQ_5 <= 1'h0;
              end else begin
                if (3'h3 == _T_1158) begin
                  portQ_5 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1158) begin
                    portQ_5 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1158) begin
                      portQ_5 <= io_bbStorePorts_1;
                    end else begin
                      portQ_5 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        if (3'h7 == _T_1176) begin
          portQ_6 <= 1'h0;
        end else begin
          if (3'h6 == _T_1176) begin
            portQ_6 <= 1'h0;
          end else begin
            if (3'h5 == _T_1176) begin
              portQ_6 <= 1'h0;
            end else begin
              if (3'h4 == _T_1176) begin
                portQ_6 <= 1'h0;
              end else begin
                if (3'h3 == _T_1176) begin
                  portQ_6 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1176) begin
                    portQ_6 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1176) begin
                      portQ_6 <= io_bbStorePorts_1;
                    end else begin
                      portQ_6 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        if (3'h7 == _T_1194) begin
          portQ_7 <= 1'h0;
        end else begin
          if (3'h6 == _T_1194) begin
            portQ_7 <= 1'h0;
          end else begin
            if (3'h5 == _T_1194) begin
              portQ_7 <= 1'h0;
            end else begin
              if (3'h4 == _T_1194) begin
                portQ_7 <= 1'h0;
              end else begin
                if (3'h3 == _T_1194) begin
                  portQ_7 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1194) begin
                    portQ_7 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1194) begin
                      portQ_7 <= io_bbStorePorts_1;
                    end else begin
                      portQ_7 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_4669) begin
          if (_T_4671) begin
            addrQ_0 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_0 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_4717) begin
          if (_T_4719) begin
            addrQ_1 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_1 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_4765) begin
          if (_T_4767) begin
            addrQ_2 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_2 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_4813) begin
          if (_T_4815) begin
            addrQ_3 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_3 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_4861) begin
          if (_T_4863) begin
            addrQ_4 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_4 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_4909) begin
          if (_T_4911) begin
            addrQ_5 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_5 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_4957) begin
          if (_T_4959) begin
            addrQ_6 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_6 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_5005) begin
          if (_T_5007) begin
            addrQ_7 <= io_addressFromStorePorts_1;
          end else begin
            addrQ_7 <= io_addressFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_4692) begin
          if (_T_4694) begin
            dataQ_0 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_0 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_4740) begin
          if (_T_4742) begin
            dataQ_1 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_1 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_4788) begin
          if (_T_4790) begin
            dataQ_2 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_2 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_4836) begin
          if (_T_4838) begin
            dataQ_3 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_3 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_4884) begin
          if (_T_4886) begin
            dataQ_4 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_4 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_4932) begin
          if (_T_4934) begin
            dataQ_5 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_5 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_4980) begin
          if (_T_4982) begin
            dataQ_6 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_6 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_5028) begin
          if (_T_5030) begin
            dataQ_7 <= io_dataFromStorePorts_1;
          end else begin
            dataQ_7 <= io_dataFromStorePorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_4669) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_4717) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_4765) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_4813) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_4861) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_4909) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_4957) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_5005) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_4692) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_4740) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_4788) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_4836) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_4884) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_4932) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_4980) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_5028) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1038;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1039;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1040;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1041;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1042;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1043;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1044;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1045;
    end
    if (reset) begin
      storeCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        storeCompleted_0 <= 1'h0;
      end else begin
        if (_T_1955) begin
          storeCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        storeCompleted_1 <= 1'h0;
      end else begin
        if (_T_1961) begin
          storeCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        storeCompleted_2 <= 1'h0;
      end else begin
        if (_T_1967) begin
          storeCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        storeCompleted_3 <= 1'h0;
      end else begin
        if (_T_1973) begin
          storeCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        storeCompleted_4 <= 1'h0;
      end else begin
        if (_T_1979) begin
          storeCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        storeCompleted_5 <= 1'h0;
      end else begin
        if (_T_1985) begin
          storeCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        storeCompleted_6 <= 1'h0;
      end else begin
        if (_T_1991) begin
          storeCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        storeCompleted_7 <= 1'h0;
      end else begin
        if (_T_1997) begin
          storeCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_1221;
      end else begin
        if (io_loadEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_1225) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_1233) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_1251;
      end else begin
        if (io_loadEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_1255) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_1263) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_1281;
      end else begin
        if (io_loadEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_1285) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_1293) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_1311;
      end else begin
        if (io_loadEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_1315) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_1323) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_1341;
      end else begin
        if (io_loadEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_1345) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_1353) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_1371;
      end else begin
        if (io_loadEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_1375) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_1383) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_1401;
      end else begin
        if (io_loadEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_1405) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_1413) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_1431;
      end else begin
        if (io_loadEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_1435) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_1443) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    previousLoadHead <= io_loadHead;
  end
endmodule
module LOAD_QUEUE_LSQ_A( // @[:@2762.2]
  input         clock, // @[:@2763.4]
  input         reset, // @[:@2764.4]
  input         io_bbStart, // @[:@2765.4]
  input  [2:0]  io_bbLoadOffsets_0, // @[:@2765.4]
  input  [2:0]  io_bbLoadOffsets_1, // @[:@2765.4]
  input  [2:0]  io_bbLoadOffsets_2, // @[:@2765.4]
  input  [2:0]  io_bbLoadOffsets_3, // @[:@2765.4]
  input  [2:0]  io_bbLoadOffsets_4, // @[:@2765.4]
  input  [2:0]  io_bbLoadOffsets_5, // @[:@2765.4]
  input  [2:0]  io_bbLoadOffsets_6, // @[:@2765.4]
  input  [2:0]  io_bbLoadOffsets_7, // @[:@2765.4]
  input         io_bbLoadPorts_1, // @[:@2765.4]
  input  [1:0]  io_bbNumLoads, // @[:@2765.4]
  output [2:0]  io_loadTail, // @[:@2765.4]
  output [2:0]  io_loadHead, // @[:@2765.4]
  output        io_loadEmpty, // @[:@2765.4]
  input  [2:0]  io_storeTail, // @[:@2765.4]
  input  [2:0]  io_storeHead, // @[:@2765.4]
  input         io_storeEmpty, // @[:@2765.4]
  input         io_storeAddrDone_0, // @[:@2765.4]
  input         io_storeAddrDone_1, // @[:@2765.4]
  input         io_storeAddrDone_2, // @[:@2765.4]
  input         io_storeAddrDone_3, // @[:@2765.4]
  input         io_storeAddrDone_4, // @[:@2765.4]
  input         io_storeAddrDone_5, // @[:@2765.4]
  input         io_storeAddrDone_6, // @[:@2765.4]
  input         io_storeAddrDone_7, // @[:@2765.4]
  input         io_storeDataDone_0, // @[:@2765.4]
  input         io_storeDataDone_1, // @[:@2765.4]
  input         io_storeDataDone_2, // @[:@2765.4]
  input         io_storeDataDone_3, // @[:@2765.4]
  input         io_storeDataDone_4, // @[:@2765.4]
  input         io_storeDataDone_5, // @[:@2765.4]
  input         io_storeDataDone_6, // @[:@2765.4]
  input         io_storeDataDone_7, // @[:@2765.4]
  input  [31:0] io_storeAddrQueue_0, // @[:@2765.4]
  input  [31:0] io_storeAddrQueue_1, // @[:@2765.4]
  input  [31:0] io_storeAddrQueue_2, // @[:@2765.4]
  input  [31:0] io_storeAddrQueue_3, // @[:@2765.4]
  input  [31:0] io_storeAddrQueue_4, // @[:@2765.4]
  input  [31:0] io_storeAddrQueue_5, // @[:@2765.4]
  input  [31:0] io_storeAddrQueue_6, // @[:@2765.4]
  input  [31:0] io_storeAddrQueue_7, // @[:@2765.4]
  input  [31:0] io_storeDataQueue_0, // @[:@2765.4]
  input  [31:0] io_storeDataQueue_1, // @[:@2765.4]
  input  [31:0] io_storeDataQueue_2, // @[:@2765.4]
  input  [31:0] io_storeDataQueue_3, // @[:@2765.4]
  input  [31:0] io_storeDataQueue_4, // @[:@2765.4]
  input  [31:0] io_storeDataQueue_5, // @[:@2765.4]
  input  [31:0] io_storeDataQueue_6, // @[:@2765.4]
  input  [31:0] io_storeDataQueue_7, // @[:@2765.4]
  output        io_loadAddrDone_0, // @[:@2765.4]
  output        io_loadAddrDone_1, // @[:@2765.4]
  output        io_loadAddrDone_2, // @[:@2765.4]
  output        io_loadAddrDone_3, // @[:@2765.4]
  output        io_loadAddrDone_4, // @[:@2765.4]
  output        io_loadAddrDone_5, // @[:@2765.4]
  output        io_loadAddrDone_6, // @[:@2765.4]
  output        io_loadAddrDone_7, // @[:@2765.4]
  output        io_loadDataDone_0, // @[:@2765.4]
  output        io_loadDataDone_1, // @[:@2765.4]
  output        io_loadDataDone_2, // @[:@2765.4]
  output        io_loadDataDone_3, // @[:@2765.4]
  output        io_loadDataDone_4, // @[:@2765.4]
  output        io_loadDataDone_5, // @[:@2765.4]
  output        io_loadDataDone_6, // @[:@2765.4]
  output        io_loadDataDone_7, // @[:@2765.4]
  output [31:0] io_loadAddrQueue_0, // @[:@2765.4]
  output [31:0] io_loadAddrQueue_1, // @[:@2765.4]
  output [31:0] io_loadAddrQueue_2, // @[:@2765.4]
  output [31:0] io_loadAddrQueue_3, // @[:@2765.4]
  output [31:0] io_loadAddrQueue_4, // @[:@2765.4]
  output [31:0] io_loadAddrQueue_5, // @[:@2765.4]
  output [31:0] io_loadAddrQueue_6, // @[:@2765.4]
  output [31:0] io_loadAddrQueue_7, // @[:@2765.4]
  input         io_loadAddrEnable_0, // @[:@2765.4]
  input         io_loadAddrEnable_1, // @[:@2765.4]
  input  [31:0] io_addrFromLoadPorts_0, // @[:@2765.4]
  input  [31:0] io_addrFromLoadPorts_1, // @[:@2765.4]
  input         io_loadPorts_0_ready, // @[:@2765.4]
  output        io_loadPorts_0_valid, // @[:@2765.4]
  output [31:0] io_loadPorts_0_bits, // @[:@2765.4]
  input         io_loadPorts_1_ready, // @[:@2765.4]
  output        io_loadPorts_1_valid, // @[:@2765.4]
  output [31:0] io_loadPorts_1_bits, // @[:@2765.4]
  input  [31:0] io_loadDataFromMem, // @[:@2765.4]
  output [31:0] io_loadAddrToMem, // @[:@2765.4]
  output        io_loadEnableToMem, // @[:@2765.4]
  input         io_memIsReadyForLoads // @[:@2765.4]
);
  reg [2:0] head; // @[LoadQueue.scala 50:21:@2767.4]
  reg [31:0] _RAND_0;
  reg [2:0] tail; // @[LoadQueue.scala 51:21:@2768.4]
  reg [31:0] _RAND_1;
  reg [2:0] offsetQ_0; // @[LoadQueue.scala 53:24:@2778.4]
  reg [31:0] _RAND_2;
  reg [2:0] offsetQ_1; // @[LoadQueue.scala 53:24:@2778.4]
  reg [31:0] _RAND_3;
  reg [2:0] offsetQ_2; // @[LoadQueue.scala 53:24:@2778.4]
  reg [31:0] _RAND_4;
  reg [2:0] offsetQ_3; // @[LoadQueue.scala 53:24:@2778.4]
  reg [31:0] _RAND_5;
  reg [2:0] offsetQ_4; // @[LoadQueue.scala 53:24:@2778.4]
  reg [31:0] _RAND_6;
  reg [2:0] offsetQ_5; // @[LoadQueue.scala 53:24:@2778.4]
  reg [31:0] _RAND_7;
  reg [2:0] offsetQ_6; // @[LoadQueue.scala 53:24:@2778.4]
  reg [31:0] _RAND_8;
  reg [2:0] offsetQ_7; // @[LoadQueue.scala 53:24:@2778.4]
  reg [31:0] _RAND_9;
  reg  portQ_0; // @[LoadQueue.scala 54:22:@2788.4]
  reg [31:0] _RAND_10;
  reg  portQ_1; // @[LoadQueue.scala 54:22:@2788.4]
  reg [31:0] _RAND_11;
  reg  portQ_2; // @[LoadQueue.scala 54:22:@2788.4]
  reg [31:0] _RAND_12;
  reg  portQ_3; // @[LoadQueue.scala 54:22:@2788.4]
  reg [31:0] _RAND_13;
  reg  portQ_4; // @[LoadQueue.scala 54:22:@2788.4]
  reg [31:0] _RAND_14;
  reg  portQ_5; // @[LoadQueue.scala 54:22:@2788.4]
  reg [31:0] _RAND_15;
  reg  portQ_6; // @[LoadQueue.scala 54:22:@2788.4]
  reg [31:0] _RAND_16;
  reg  portQ_7; // @[LoadQueue.scala 54:22:@2788.4]
  reg [31:0] _RAND_17;
  reg [31:0] addrQ_0; // @[LoadQueue.scala 55:22:@2798.4]
  reg [31:0] _RAND_18;
  reg [31:0] addrQ_1; // @[LoadQueue.scala 55:22:@2798.4]
  reg [31:0] _RAND_19;
  reg [31:0] addrQ_2; // @[LoadQueue.scala 55:22:@2798.4]
  reg [31:0] _RAND_20;
  reg [31:0] addrQ_3; // @[LoadQueue.scala 55:22:@2798.4]
  reg [31:0] _RAND_21;
  reg [31:0] addrQ_4; // @[LoadQueue.scala 55:22:@2798.4]
  reg [31:0] _RAND_22;
  reg [31:0] addrQ_5; // @[LoadQueue.scala 55:22:@2798.4]
  reg [31:0] _RAND_23;
  reg [31:0] addrQ_6; // @[LoadQueue.scala 55:22:@2798.4]
  reg [31:0] _RAND_24;
  reg [31:0] addrQ_7; // @[LoadQueue.scala 55:22:@2798.4]
  reg [31:0] _RAND_25;
  reg [31:0] dataQ_0; // @[LoadQueue.scala 56:22:@2808.4]
  reg [31:0] _RAND_26;
  reg [31:0] dataQ_1; // @[LoadQueue.scala 56:22:@2808.4]
  reg [31:0] _RAND_27;
  reg [31:0] dataQ_2; // @[LoadQueue.scala 56:22:@2808.4]
  reg [31:0] _RAND_28;
  reg [31:0] dataQ_3; // @[LoadQueue.scala 56:22:@2808.4]
  reg [31:0] _RAND_29;
  reg [31:0] dataQ_4; // @[LoadQueue.scala 56:22:@2808.4]
  reg [31:0] _RAND_30;
  reg [31:0] dataQ_5; // @[LoadQueue.scala 56:22:@2808.4]
  reg [31:0] _RAND_31;
  reg [31:0] dataQ_6; // @[LoadQueue.scala 56:22:@2808.4]
  reg [31:0] _RAND_32;
  reg [31:0] dataQ_7; // @[LoadQueue.scala 56:22:@2808.4]
  reg [31:0] _RAND_33;
  reg  addrKnown_0; // @[LoadQueue.scala 57:26:@2818.4]
  reg [31:0] _RAND_34;
  reg  addrKnown_1; // @[LoadQueue.scala 57:26:@2818.4]
  reg [31:0] _RAND_35;
  reg  addrKnown_2; // @[LoadQueue.scala 57:26:@2818.4]
  reg [31:0] _RAND_36;
  reg  addrKnown_3; // @[LoadQueue.scala 57:26:@2818.4]
  reg [31:0] _RAND_37;
  reg  addrKnown_4; // @[LoadQueue.scala 57:26:@2818.4]
  reg [31:0] _RAND_38;
  reg  addrKnown_5; // @[LoadQueue.scala 57:26:@2818.4]
  reg [31:0] _RAND_39;
  reg  addrKnown_6; // @[LoadQueue.scala 57:26:@2818.4]
  reg [31:0] _RAND_40;
  reg  addrKnown_7; // @[LoadQueue.scala 57:26:@2818.4]
  reg [31:0] _RAND_41;
  reg  dataKnown_0; // @[LoadQueue.scala 58:26:@2828.4]
  reg [31:0] _RAND_42;
  reg  dataKnown_1; // @[LoadQueue.scala 58:26:@2828.4]
  reg [31:0] _RAND_43;
  reg  dataKnown_2; // @[LoadQueue.scala 58:26:@2828.4]
  reg [31:0] _RAND_44;
  reg  dataKnown_3; // @[LoadQueue.scala 58:26:@2828.4]
  reg [31:0] _RAND_45;
  reg  dataKnown_4; // @[LoadQueue.scala 58:26:@2828.4]
  reg [31:0] _RAND_46;
  reg  dataKnown_5; // @[LoadQueue.scala 58:26:@2828.4]
  reg [31:0] _RAND_47;
  reg  dataKnown_6; // @[LoadQueue.scala 58:26:@2828.4]
  reg [31:0] _RAND_48;
  reg  dataKnown_7; // @[LoadQueue.scala 58:26:@2828.4]
  reg [31:0] _RAND_49;
  reg  loadCompleted_0; // @[LoadQueue.scala 59:30:@2838.4]
  reg [31:0] _RAND_50;
  reg  loadCompleted_1; // @[LoadQueue.scala 59:30:@2838.4]
  reg [31:0] _RAND_51;
  reg  loadCompleted_2; // @[LoadQueue.scala 59:30:@2838.4]
  reg [31:0] _RAND_52;
  reg  loadCompleted_3; // @[LoadQueue.scala 59:30:@2838.4]
  reg [31:0] _RAND_53;
  reg  loadCompleted_4; // @[LoadQueue.scala 59:30:@2838.4]
  reg [31:0] _RAND_54;
  reg  loadCompleted_5; // @[LoadQueue.scala 59:30:@2838.4]
  reg [31:0] _RAND_55;
  reg  loadCompleted_6; // @[LoadQueue.scala 59:30:@2838.4]
  reg [31:0] _RAND_56;
  reg  loadCompleted_7; // @[LoadQueue.scala 59:30:@2838.4]
  reg [31:0] _RAND_57;
  reg  allocatedEntries_0; // @[LoadQueue.scala 60:33:@2848.4]
  reg [31:0] _RAND_58;
  reg  allocatedEntries_1; // @[LoadQueue.scala 60:33:@2848.4]
  reg [31:0] _RAND_59;
  reg  allocatedEntries_2; // @[LoadQueue.scala 60:33:@2848.4]
  reg [31:0] _RAND_60;
  reg  allocatedEntries_3; // @[LoadQueue.scala 60:33:@2848.4]
  reg [31:0] _RAND_61;
  reg  allocatedEntries_4; // @[LoadQueue.scala 60:33:@2848.4]
  reg [31:0] _RAND_62;
  reg  allocatedEntries_5; // @[LoadQueue.scala 60:33:@2848.4]
  reg [31:0] _RAND_63;
  reg  allocatedEntries_6; // @[LoadQueue.scala 60:33:@2848.4]
  reg [31:0] _RAND_64;
  reg  allocatedEntries_7; // @[LoadQueue.scala 60:33:@2848.4]
  reg [31:0] _RAND_65;
  reg  bypassInitiated_0; // @[LoadQueue.scala 61:32:@2858.4]
  reg [31:0] _RAND_66;
  reg  bypassInitiated_1; // @[LoadQueue.scala 61:32:@2858.4]
  reg [31:0] _RAND_67;
  reg  bypassInitiated_2; // @[LoadQueue.scala 61:32:@2858.4]
  reg [31:0] _RAND_68;
  reg  bypassInitiated_3; // @[LoadQueue.scala 61:32:@2858.4]
  reg [31:0] _RAND_69;
  reg  bypassInitiated_4; // @[LoadQueue.scala 61:32:@2858.4]
  reg [31:0] _RAND_70;
  reg  bypassInitiated_5; // @[LoadQueue.scala 61:32:@2858.4]
  reg [31:0] _RAND_71;
  reg  bypassInitiated_6; // @[LoadQueue.scala 61:32:@2858.4]
  reg [31:0] _RAND_72;
  reg  bypassInitiated_7; // @[LoadQueue.scala 61:32:@2858.4]
  reg [31:0] _RAND_73;
  reg  checkBits_0; // @[LoadQueue.scala 62:26:@2868.4]
  reg [31:0] _RAND_74;
  reg  checkBits_1; // @[LoadQueue.scala 62:26:@2868.4]
  reg [31:0] _RAND_75;
  reg  checkBits_2; // @[LoadQueue.scala 62:26:@2868.4]
  reg [31:0] _RAND_76;
  reg  checkBits_3; // @[LoadQueue.scala 62:26:@2868.4]
  reg [31:0] _RAND_77;
  reg  checkBits_4; // @[LoadQueue.scala 62:26:@2868.4]
  reg [31:0] _RAND_78;
  reg  checkBits_5; // @[LoadQueue.scala 62:26:@2868.4]
  reg [31:0] _RAND_79;
  reg  checkBits_6; // @[LoadQueue.scala 62:26:@2868.4]
  reg [31:0] _RAND_80;
  reg  checkBits_7; // @[LoadQueue.scala 62:26:@2868.4]
  reg [31:0] _RAND_81;
  wire [4:0] _GEN_712; // @[util.scala 14:20:@2870.4]
  wire [5:0] _T_1020; // @[util.scala 14:20:@2870.4]
  wire [5:0] _T_1021; // @[util.scala 14:20:@2871.4]
  wire [4:0] _T_1022; // @[util.scala 14:20:@2872.4]
  wire [4:0] _GEN_0; // @[util.scala 14:25:@2873.4]
  wire [3:0] _T_1023; // @[util.scala 14:25:@2873.4]
  wire [3:0] _GEN_713; // @[LoadQueue.scala 71:46:@2874.4]
  wire  _T_1024; // @[LoadQueue.scala 71:46:@2874.4]
  wire  initBits_0; // @[LoadQueue.scala 71:63:@2875.4]
  wire [5:0] _T_1029; // @[util.scala 14:20:@2877.4]
  wire [5:0] _T_1030; // @[util.scala 14:20:@2878.4]
  wire [4:0] _T_1031; // @[util.scala 14:20:@2879.4]
  wire [4:0] _GEN_8; // @[util.scala 14:25:@2880.4]
  wire [3:0] _T_1032; // @[util.scala 14:25:@2880.4]
  wire  _T_1033; // @[LoadQueue.scala 71:46:@2881.4]
  wire  initBits_1; // @[LoadQueue.scala 71:63:@2882.4]
  wire [5:0] _T_1038; // @[util.scala 14:20:@2884.4]
  wire [5:0] _T_1039; // @[util.scala 14:20:@2885.4]
  wire [4:0] _T_1040; // @[util.scala 14:20:@2886.4]
  wire [4:0] _GEN_18; // @[util.scala 14:25:@2887.4]
  wire [3:0] _T_1041; // @[util.scala 14:25:@2887.4]
  wire  _T_1042; // @[LoadQueue.scala 71:46:@2888.4]
  wire  initBits_2; // @[LoadQueue.scala 71:63:@2889.4]
  wire [5:0] _T_1047; // @[util.scala 14:20:@2891.4]
  wire [5:0] _T_1048; // @[util.scala 14:20:@2892.4]
  wire [4:0] _T_1049; // @[util.scala 14:20:@2893.4]
  wire [4:0] _GEN_26; // @[util.scala 14:25:@2894.4]
  wire [3:0] _T_1050; // @[util.scala 14:25:@2894.4]
  wire  _T_1051; // @[LoadQueue.scala 71:46:@2895.4]
  wire  initBits_3; // @[LoadQueue.scala 71:63:@2896.4]
  wire [5:0] _T_1056; // @[util.scala 14:20:@2898.4]
  wire [5:0] _T_1057; // @[util.scala 14:20:@2899.4]
  wire [4:0] _T_1058; // @[util.scala 14:20:@2900.4]
  wire [4:0] _GEN_36; // @[util.scala 14:25:@2901.4]
  wire [3:0] _T_1059; // @[util.scala 14:25:@2901.4]
  wire  _T_1060; // @[LoadQueue.scala 71:46:@2902.4]
  wire  initBits_4; // @[LoadQueue.scala 71:63:@2903.4]
  wire [5:0] _T_1065; // @[util.scala 14:20:@2905.4]
  wire [5:0] _T_1066; // @[util.scala 14:20:@2906.4]
  wire [4:0] _T_1067; // @[util.scala 14:20:@2907.4]
  wire [4:0] _GEN_44; // @[util.scala 14:25:@2908.4]
  wire [3:0] _T_1068; // @[util.scala 14:25:@2908.4]
  wire  _T_1069; // @[LoadQueue.scala 71:46:@2909.4]
  wire  initBits_5; // @[LoadQueue.scala 71:63:@2910.4]
  wire [5:0] _T_1074; // @[util.scala 14:20:@2912.4]
  wire [5:0] _T_1075; // @[util.scala 14:20:@2913.4]
  wire [4:0] _T_1076; // @[util.scala 14:20:@2914.4]
  wire [4:0] _GEN_54; // @[util.scala 14:25:@2915.4]
  wire [3:0] _T_1077; // @[util.scala 14:25:@2915.4]
  wire  _T_1078; // @[LoadQueue.scala 71:46:@2916.4]
  wire  initBits_6; // @[LoadQueue.scala 71:63:@2917.4]
  wire [5:0] _T_1083; // @[util.scala 14:20:@2919.4]
  wire [5:0] _T_1084; // @[util.scala 14:20:@2920.4]
  wire [4:0] _T_1085; // @[util.scala 14:20:@2921.4]
  wire [4:0] _GEN_62; // @[util.scala 14:25:@2922.4]
  wire [3:0] _T_1086; // @[util.scala 14:25:@2922.4]
  wire  _T_1087; // @[LoadQueue.scala 71:46:@2923.4]
  wire  initBits_7; // @[LoadQueue.scala 71:63:@2924.4]
  wire  _T_1102; // @[LoadQueue.scala 73:78:@2934.4]
  wire  _T_1103; // @[LoadQueue.scala 73:78:@2935.4]
  wire  _T_1104; // @[LoadQueue.scala 73:78:@2936.4]
  wire  _T_1105; // @[LoadQueue.scala 73:78:@2937.4]
  wire  _T_1106; // @[LoadQueue.scala 73:78:@2938.4]
  wire  _T_1107; // @[LoadQueue.scala 73:78:@2939.4]
  wire  _T_1108; // @[LoadQueue.scala 73:78:@2940.4]
  wire  _T_1109; // @[LoadQueue.scala 73:78:@2941.4]
  wire [2:0] _T_1132; // @[:@2965.6]
  wire [2:0] _GEN_1; // @[LoadQueue.scala 77:20:@2966.6]
  wire [2:0] _GEN_2; // @[LoadQueue.scala 77:20:@2966.6]
  wire [2:0] _GEN_3; // @[LoadQueue.scala 77:20:@2966.6]
  wire [2:0] _GEN_4; // @[LoadQueue.scala 77:20:@2966.6]
  wire [2:0] _GEN_5; // @[LoadQueue.scala 77:20:@2966.6]
  wire [2:0] _GEN_6; // @[LoadQueue.scala 77:20:@2966.6]
  wire [2:0] _GEN_7; // @[LoadQueue.scala 77:20:@2966.6]
  wire  _GEN_9; // @[LoadQueue.scala 78:18:@2973.6]
  wire  _GEN_10; // @[LoadQueue.scala 78:18:@2973.6]
  wire  _GEN_11; // @[LoadQueue.scala 78:18:@2973.6]
  wire  _GEN_12; // @[LoadQueue.scala 78:18:@2973.6]
  wire  _GEN_13; // @[LoadQueue.scala 78:18:@2973.6]
  wire  _GEN_14; // @[LoadQueue.scala 78:18:@2973.6]
  wire  _GEN_15; // @[LoadQueue.scala 78:18:@2973.6]
  wire [2:0] _GEN_16; // @[LoadQueue.scala 76:25:@2959.4]
  wire  _GEN_17; // @[LoadQueue.scala 76:25:@2959.4]
  wire [2:0] _T_1150; // @[:@2981.6]
  wire [2:0] _GEN_19; // @[LoadQueue.scala 77:20:@2982.6]
  wire [2:0] _GEN_20; // @[LoadQueue.scala 77:20:@2982.6]
  wire [2:0] _GEN_21; // @[LoadQueue.scala 77:20:@2982.6]
  wire [2:0] _GEN_22; // @[LoadQueue.scala 77:20:@2982.6]
  wire [2:0] _GEN_23; // @[LoadQueue.scala 77:20:@2982.6]
  wire [2:0] _GEN_24; // @[LoadQueue.scala 77:20:@2982.6]
  wire [2:0] _GEN_25; // @[LoadQueue.scala 77:20:@2982.6]
  wire  _GEN_27; // @[LoadQueue.scala 78:18:@2989.6]
  wire  _GEN_28; // @[LoadQueue.scala 78:18:@2989.6]
  wire  _GEN_29; // @[LoadQueue.scala 78:18:@2989.6]
  wire  _GEN_30; // @[LoadQueue.scala 78:18:@2989.6]
  wire  _GEN_31; // @[LoadQueue.scala 78:18:@2989.6]
  wire  _GEN_32; // @[LoadQueue.scala 78:18:@2989.6]
  wire  _GEN_33; // @[LoadQueue.scala 78:18:@2989.6]
  wire [2:0] _GEN_34; // @[LoadQueue.scala 76:25:@2975.4]
  wire  _GEN_35; // @[LoadQueue.scala 76:25:@2975.4]
  wire [2:0] _T_1168; // @[:@2997.6]
  wire [2:0] _GEN_37; // @[LoadQueue.scala 77:20:@2998.6]
  wire [2:0] _GEN_38; // @[LoadQueue.scala 77:20:@2998.6]
  wire [2:0] _GEN_39; // @[LoadQueue.scala 77:20:@2998.6]
  wire [2:0] _GEN_40; // @[LoadQueue.scala 77:20:@2998.6]
  wire [2:0] _GEN_41; // @[LoadQueue.scala 77:20:@2998.6]
  wire [2:0] _GEN_42; // @[LoadQueue.scala 77:20:@2998.6]
  wire [2:0] _GEN_43; // @[LoadQueue.scala 77:20:@2998.6]
  wire  _GEN_45; // @[LoadQueue.scala 78:18:@3005.6]
  wire  _GEN_46; // @[LoadQueue.scala 78:18:@3005.6]
  wire  _GEN_47; // @[LoadQueue.scala 78:18:@3005.6]
  wire  _GEN_48; // @[LoadQueue.scala 78:18:@3005.6]
  wire  _GEN_49; // @[LoadQueue.scala 78:18:@3005.6]
  wire  _GEN_50; // @[LoadQueue.scala 78:18:@3005.6]
  wire  _GEN_51; // @[LoadQueue.scala 78:18:@3005.6]
  wire [2:0] _GEN_52; // @[LoadQueue.scala 76:25:@2991.4]
  wire  _GEN_53; // @[LoadQueue.scala 76:25:@2991.4]
  wire [2:0] _T_1186; // @[:@3013.6]
  wire [2:0] _GEN_55; // @[LoadQueue.scala 77:20:@3014.6]
  wire [2:0] _GEN_56; // @[LoadQueue.scala 77:20:@3014.6]
  wire [2:0] _GEN_57; // @[LoadQueue.scala 77:20:@3014.6]
  wire [2:0] _GEN_58; // @[LoadQueue.scala 77:20:@3014.6]
  wire [2:0] _GEN_59; // @[LoadQueue.scala 77:20:@3014.6]
  wire [2:0] _GEN_60; // @[LoadQueue.scala 77:20:@3014.6]
  wire [2:0] _GEN_61; // @[LoadQueue.scala 77:20:@3014.6]
  wire  _GEN_63; // @[LoadQueue.scala 78:18:@3021.6]
  wire  _GEN_64; // @[LoadQueue.scala 78:18:@3021.6]
  wire  _GEN_65; // @[LoadQueue.scala 78:18:@3021.6]
  wire  _GEN_66; // @[LoadQueue.scala 78:18:@3021.6]
  wire  _GEN_67; // @[LoadQueue.scala 78:18:@3021.6]
  wire  _GEN_68; // @[LoadQueue.scala 78:18:@3021.6]
  wire  _GEN_69; // @[LoadQueue.scala 78:18:@3021.6]
  wire [2:0] _GEN_70; // @[LoadQueue.scala 76:25:@3007.4]
  wire  _GEN_71; // @[LoadQueue.scala 76:25:@3007.4]
  wire [2:0] _T_1204; // @[:@3029.6]
  wire [2:0] _GEN_73; // @[LoadQueue.scala 77:20:@3030.6]
  wire [2:0] _GEN_74; // @[LoadQueue.scala 77:20:@3030.6]
  wire [2:0] _GEN_75; // @[LoadQueue.scala 77:20:@3030.6]
  wire [2:0] _GEN_76; // @[LoadQueue.scala 77:20:@3030.6]
  wire [2:0] _GEN_77; // @[LoadQueue.scala 77:20:@3030.6]
  wire [2:0] _GEN_78; // @[LoadQueue.scala 77:20:@3030.6]
  wire [2:0] _GEN_79; // @[LoadQueue.scala 77:20:@3030.6]
  wire  _GEN_81; // @[LoadQueue.scala 78:18:@3037.6]
  wire  _GEN_82; // @[LoadQueue.scala 78:18:@3037.6]
  wire  _GEN_83; // @[LoadQueue.scala 78:18:@3037.6]
  wire  _GEN_84; // @[LoadQueue.scala 78:18:@3037.6]
  wire  _GEN_85; // @[LoadQueue.scala 78:18:@3037.6]
  wire  _GEN_86; // @[LoadQueue.scala 78:18:@3037.6]
  wire  _GEN_87; // @[LoadQueue.scala 78:18:@3037.6]
  wire [2:0] _GEN_88; // @[LoadQueue.scala 76:25:@3023.4]
  wire  _GEN_89; // @[LoadQueue.scala 76:25:@3023.4]
  wire [2:0] _T_1222; // @[:@3045.6]
  wire [2:0] _GEN_91; // @[LoadQueue.scala 77:20:@3046.6]
  wire [2:0] _GEN_92; // @[LoadQueue.scala 77:20:@3046.6]
  wire [2:0] _GEN_93; // @[LoadQueue.scala 77:20:@3046.6]
  wire [2:0] _GEN_94; // @[LoadQueue.scala 77:20:@3046.6]
  wire [2:0] _GEN_95; // @[LoadQueue.scala 77:20:@3046.6]
  wire [2:0] _GEN_96; // @[LoadQueue.scala 77:20:@3046.6]
  wire [2:0] _GEN_97; // @[LoadQueue.scala 77:20:@3046.6]
  wire  _GEN_99; // @[LoadQueue.scala 78:18:@3053.6]
  wire  _GEN_100; // @[LoadQueue.scala 78:18:@3053.6]
  wire  _GEN_101; // @[LoadQueue.scala 78:18:@3053.6]
  wire  _GEN_102; // @[LoadQueue.scala 78:18:@3053.6]
  wire  _GEN_103; // @[LoadQueue.scala 78:18:@3053.6]
  wire  _GEN_104; // @[LoadQueue.scala 78:18:@3053.6]
  wire  _GEN_105; // @[LoadQueue.scala 78:18:@3053.6]
  wire [2:0] _GEN_106; // @[LoadQueue.scala 76:25:@3039.4]
  wire  _GEN_107; // @[LoadQueue.scala 76:25:@3039.4]
  wire [2:0] _T_1240; // @[:@3061.6]
  wire [2:0] _GEN_109; // @[LoadQueue.scala 77:20:@3062.6]
  wire [2:0] _GEN_110; // @[LoadQueue.scala 77:20:@3062.6]
  wire [2:0] _GEN_111; // @[LoadQueue.scala 77:20:@3062.6]
  wire [2:0] _GEN_112; // @[LoadQueue.scala 77:20:@3062.6]
  wire [2:0] _GEN_113; // @[LoadQueue.scala 77:20:@3062.6]
  wire [2:0] _GEN_114; // @[LoadQueue.scala 77:20:@3062.6]
  wire [2:0] _GEN_115; // @[LoadQueue.scala 77:20:@3062.6]
  wire  _GEN_117; // @[LoadQueue.scala 78:18:@3069.6]
  wire  _GEN_118; // @[LoadQueue.scala 78:18:@3069.6]
  wire  _GEN_119; // @[LoadQueue.scala 78:18:@3069.6]
  wire  _GEN_120; // @[LoadQueue.scala 78:18:@3069.6]
  wire  _GEN_121; // @[LoadQueue.scala 78:18:@3069.6]
  wire  _GEN_122; // @[LoadQueue.scala 78:18:@3069.6]
  wire  _GEN_123; // @[LoadQueue.scala 78:18:@3069.6]
  wire [2:0] _GEN_124; // @[LoadQueue.scala 76:25:@3055.4]
  wire  _GEN_125; // @[LoadQueue.scala 76:25:@3055.4]
  wire [2:0] _T_1258; // @[:@3077.6]
  wire [2:0] _GEN_127; // @[LoadQueue.scala 77:20:@3078.6]
  wire [2:0] _GEN_128; // @[LoadQueue.scala 77:20:@3078.6]
  wire [2:0] _GEN_129; // @[LoadQueue.scala 77:20:@3078.6]
  wire [2:0] _GEN_130; // @[LoadQueue.scala 77:20:@3078.6]
  wire [2:0] _GEN_131; // @[LoadQueue.scala 77:20:@3078.6]
  wire [2:0] _GEN_132; // @[LoadQueue.scala 77:20:@3078.6]
  wire [2:0] _GEN_133; // @[LoadQueue.scala 77:20:@3078.6]
  wire  _GEN_135; // @[LoadQueue.scala 78:18:@3085.6]
  wire  _GEN_136; // @[LoadQueue.scala 78:18:@3085.6]
  wire  _GEN_137; // @[LoadQueue.scala 78:18:@3085.6]
  wire  _GEN_138; // @[LoadQueue.scala 78:18:@3085.6]
  wire  _GEN_139; // @[LoadQueue.scala 78:18:@3085.6]
  wire  _GEN_140; // @[LoadQueue.scala 78:18:@3085.6]
  wire  _GEN_141; // @[LoadQueue.scala 78:18:@3085.6]
  wire [2:0] _GEN_142; // @[LoadQueue.scala 76:25:@3071.4]
  wire  _GEN_143; // @[LoadQueue.scala 76:25:@3071.4]
  reg [2:0] previousStoreHead; // @[LoadQueue.scala 93:34:@3087.4]
  reg [31:0] _RAND_82;
  wire [3:0] _T_1280; // @[util.scala 10:8:@3096.6]
  wire [3:0] _GEN_72; // @[util.scala 10:14:@3097.6]
  wire [3:0] _T_1281; // @[util.scala 10:14:@3097.6]
  wire [3:0] _GEN_745; // @[LoadQueue.scala 97:56:@3098.6]
  wire  _T_1282; // @[LoadQueue.scala 97:56:@3098.6]
  wire  _T_1283; // @[LoadQueue.scala 96:50:@3099.6]
  wire  _T_1285; // @[LoadQueue.scala 96:34:@3100.6]
  wire  _T_1287; // @[LoadQueue.scala 101:36:@3108.8]
  wire  _T_1288; // @[LoadQueue.scala 101:86:@3109.8]
  wire  _T_1289; // @[LoadQueue.scala 101:61:@3110.8]
  wire  _T_1291; // @[LoadQueue.scala 103:36:@3115.10]
  wire  _T_1292; // @[LoadQueue.scala 103:69:@3116.10]
  wire  _T_1293; // @[LoadQueue.scala 104:31:@3117.10]
  wire  _T_1294; // @[LoadQueue.scala 103:94:@3118.10]
  wire  _T_1296; // @[LoadQueue.scala 103:54:@3119.10]
  wire  _T_1297; // @[LoadQueue.scala 103:51:@3120.10]
  wire  _GEN_152; // @[LoadQueue.scala 104:53:@3121.10]
  wire  _GEN_153; // @[LoadQueue.scala 101:102:@3111.8]
  wire  _GEN_154; // @[LoadQueue.scala 99:27:@3104.6]
  wire  _GEN_155; // @[LoadQueue.scala 95:34:@3089.4]
  wire [3:0] _T_1310; // @[util.scala 10:8:@3132.6]
  wire [3:0] _GEN_80; // @[util.scala 10:14:@3133.6]
  wire [3:0] _T_1311; // @[util.scala 10:14:@3133.6]
  wire  _T_1312; // @[LoadQueue.scala 97:56:@3134.6]
  wire  _T_1313; // @[LoadQueue.scala 96:50:@3135.6]
  wire  _T_1315; // @[LoadQueue.scala 96:34:@3136.6]
  wire  _T_1317; // @[LoadQueue.scala 101:36:@3144.8]
  wire  _T_1318; // @[LoadQueue.scala 101:86:@3145.8]
  wire  _T_1319; // @[LoadQueue.scala 101:61:@3146.8]
  wire  _T_1322; // @[LoadQueue.scala 103:69:@3152.10]
  wire  _T_1323; // @[LoadQueue.scala 104:31:@3153.10]
  wire  _T_1324; // @[LoadQueue.scala 103:94:@3154.10]
  wire  _T_1326; // @[LoadQueue.scala 103:54:@3155.10]
  wire  _T_1327; // @[LoadQueue.scala 103:51:@3156.10]
  wire  _GEN_164; // @[LoadQueue.scala 104:53:@3157.10]
  wire  _GEN_165; // @[LoadQueue.scala 101:102:@3147.8]
  wire  _GEN_166; // @[LoadQueue.scala 99:27:@3140.6]
  wire  _GEN_167; // @[LoadQueue.scala 95:34:@3125.4]
  wire [3:0] _T_1340; // @[util.scala 10:8:@3168.6]
  wire [3:0] _GEN_90; // @[util.scala 10:14:@3169.6]
  wire [3:0] _T_1341; // @[util.scala 10:14:@3169.6]
  wire  _T_1342; // @[LoadQueue.scala 97:56:@3170.6]
  wire  _T_1343; // @[LoadQueue.scala 96:50:@3171.6]
  wire  _T_1345; // @[LoadQueue.scala 96:34:@3172.6]
  wire  _T_1347; // @[LoadQueue.scala 101:36:@3180.8]
  wire  _T_1348; // @[LoadQueue.scala 101:86:@3181.8]
  wire  _T_1349; // @[LoadQueue.scala 101:61:@3182.8]
  wire  _T_1352; // @[LoadQueue.scala 103:69:@3188.10]
  wire  _T_1353; // @[LoadQueue.scala 104:31:@3189.10]
  wire  _T_1354; // @[LoadQueue.scala 103:94:@3190.10]
  wire  _T_1356; // @[LoadQueue.scala 103:54:@3191.10]
  wire  _T_1357; // @[LoadQueue.scala 103:51:@3192.10]
  wire  _GEN_176; // @[LoadQueue.scala 104:53:@3193.10]
  wire  _GEN_177; // @[LoadQueue.scala 101:102:@3183.8]
  wire  _GEN_178; // @[LoadQueue.scala 99:27:@3176.6]
  wire  _GEN_179; // @[LoadQueue.scala 95:34:@3161.4]
  wire [3:0] _T_1370; // @[util.scala 10:8:@3204.6]
  wire [3:0] _GEN_98; // @[util.scala 10:14:@3205.6]
  wire [3:0] _T_1371; // @[util.scala 10:14:@3205.6]
  wire  _T_1372; // @[LoadQueue.scala 97:56:@3206.6]
  wire  _T_1373; // @[LoadQueue.scala 96:50:@3207.6]
  wire  _T_1375; // @[LoadQueue.scala 96:34:@3208.6]
  wire  _T_1377; // @[LoadQueue.scala 101:36:@3216.8]
  wire  _T_1378; // @[LoadQueue.scala 101:86:@3217.8]
  wire  _T_1379; // @[LoadQueue.scala 101:61:@3218.8]
  wire  _T_1382; // @[LoadQueue.scala 103:69:@3224.10]
  wire  _T_1383; // @[LoadQueue.scala 104:31:@3225.10]
  wire  _T_1384; // @[LoadQueue.scala 103:94:@3226.10]
  wire  _T_1386; // @[LoadQueue.scala 103:54:@3227.10]
  wire  _T_1387; // @[LoadQueue.scala 103:51:@3228.10]
  wire  _GEN_188; // @[LoadQueue.scala 104:53:@3229.10]
  wire  _GEN_189; // @[LoadQueue.scala 101:102:@3219.8]
  wire  _GEN_190; // @[LoadQueue.scala 99:27:@3212.6]
  wire  _GEN_191; // @[LoadQueue.scala 95:34:@3197.4]
  wire [3:0] _T_1400; // @[util.scala 10:8:@3240.6]
  wire [3:0] _GEN_108; // @[util.scala 10:14:@3241.6]
  wire [3:0] _T_1401; // @[util.scala 10:14:@3241.6]
  wire  _T_1402; // @[LoadQueue.scala 97:56:@3242.6]
  wire  _T_1403; // @[LoadQueue.scala 96:50:@3243.6]
  wire  _T_1405; // @[LoadQueue.scala 96:34:@3244.6]
  wire  _T_1407; // @[LoadQueue.scala 101:36:@3252.8]
  wire  _T_1408; // @[LoadQueue.scala 101:86:@3253.8]
  wire  _T_1409; // @[LoadQueue.scala 101:61:@3254.8]
  wire  _T_1412; // @[LoadQueue.scala 103:69:@3260.10]
  wire  _T_1413; // @[LoadQueue.scala 104:31:@3261.10]
  wire  _T_1414; // @[LoadQueue.scala 103:94:@3262.10]
  wire  _T_1416; // @[LoadQueue.scala 103:54:@3263.10]
  wire  _T_1417; // @[LoadQueue.scala 103:51:@3264.10]
  wire  _GEN_200; // @[LoadQueue.scala 104:53:@3265.10]
  wire  _GEN_201; // @[LoadQueue.scala 101:102:@3255.8]
  wire  _GEN_202; // @[LoadQueue.scala 99:27:@3248.6]
  wire  _GEN_203; // @[LoadQueue.scala 95:34:@3233.4]
  wire [3:0] _T_1430; // @[util.scala 10:8:@3276.6]
  wire [3:0] _GEN_116; // @[util.scala 10:14:@3277.6]
  wire [3:0] _T_1431; // @[util.scala 10:14:@3277.6]
  wire  _T_1432; // @[LoadQueue.scala 97:56:@3278.6]
  wire  _T_1433; // @[LoadQueue.scala 96:50:@3279.6]
  wire  _T_1435; // @[LoadQueue.scala 96:34:@3280.6]
  wire  _T_1437; // @[LoadQueue.scala 101:36:@3288.8]
  wire  _T_1438; // @[LoadQueue.scala 101:86:@3289.8]
  wire  _T_1439; // @[LoadQueue.scala 101:61:@3290.8]
  wire  _T_1442; // @[LoadQueue.scala 103:69:@3296.10]
  wire  _T_1443; // @[LoadQueue.scala 104:31:@3297.10]
  wire  _T_1444; // @[LoadQueue.scala 103:94:@3298.10]
  wire  _T_1446; // @[LoadQueue.scala 103:54:@3299.10]
  wire  _T_1447; // @[LoadQueue.scala 103:51:@3300.10]
  wire  _GEN_212; // @[LoadQueue.scala 104:53:@3301.10]
  wire  _GEN_213; // @[LoadQueue.scala 101:102:@3291.8]
  wire  _GEN_214; // @[LoadQueue.scala 99:27:@3284.6]
  wire  _GEN_215; // @[LoadQueue.scala 95:34:@3269.4]
  wire [3:0] _T_1460; // @[util.scala 10:8:@3312.6]
  wire [3:0] _GEN_126; // @[util.scala 10:14:@3313.6]
  wire [3:0] _T_1461; // @[util.scala 10:14:@3313.6]
  wire  _T_1462; // @[LoadQueue.scala 97:56:@3314.6]
  wire  _T_1463; // @[LoadQueue.scala 96:50:@3315.6]
  wire  _T_1465; // @[LoadQueue.scala 96:34:@3316.6]
  wire  _T_1467; // @[LoadQueue.scala 101:36:@3324.8]
  wire  _T_1468; // @[LoadQueue.scala 101:86:@3325.8]
  wire  _T_1469; // @[LoadQueue.scala 101:61:@3326.8]
  wire  _T_1472; // @[LoadQueue.scala 103:69:@3332.10]
  wire  _T_1473; // @[LoadQueue.scala 104:31:@3333.10]
  wire  _T_1474; // @[LoadQueue.scala 103:94:@3334.10]
  wire  _T_1476; // @[LoadQueue.scala 103:54:@3335.10]
  wire  _T_1477; // @[LoadQueue.scala 103:51:@3336.10]
  wire  _GEN_224; // @[LoadQueue.scala 104:53:@3337.10]
  wire  _GEN_225; // @[LoadQueue.scala 101:102:@3327.8]
  wire  _GEN_226; // @[LoadQueue.scala 99:27:@3320.6]
  wire  _GEN_227; // @[LoadQueue.scala 95:34:@3305.4]
  wire [3:0] _T_1490; // @[util.scala 10:8:@3348.6]
  wire [3:0] _GEN_134; // @[util.scala 10:14:@3349.6]
  wire [3:0] _T_1491; // @[util.scala 10:14:@3349.6]
  wire  _T_1492; // @[LoadQueue.scala 97:56:@3350.6]
  wire  _T_1493; // @[LoadQueue.scala 96:50:@3351.6]
  wire  _T_1495; // @[LoadQueue.scala 96:34:@3352.6]
  wire  _T_1497; // @[LoadQueue.scala 101:36:@3360.8]
  wire  _T_1498; // @[LoadQueue.scala 101:86:@3361.8]
  wire  _T_1499; // @[LoadQueue.scala 101:61:@3362.8]
  wire  _T_1502; // @[LoadQueue.scala 103:69:@3368.10]
  wire  _T_1503; // @[LoadQueue.scala 104:31:@3369.10]
  wire  _T_1504; // @[LoadQueue.scala 103:94:@3370.10]
  wire  _T_1506; // @[LoadQueue.scala 103:54:@3371.10]
  wire  _T_1507; // @[LoadQueue.scala 103:51:@3372.10]
  wire  _GEN_236; // @[LoadQueue.scala 104:53:@3373.10]
  wire  _GEN_237; // @[LoadQueue.scala 101:102:@3363.8]
  wire  _GEN_238; // @[LoadQueue.scala 99:27:@3356.6]
  wire  _GEN_239; // @[LoadQueue.scala 95:34:@3341.4]
  wire [7:0] _T_1511; // @[OneHot.scala 52:12:@3378.4]
  wire  _T_1513; // @[util.scala 60:60:@3380.4]
  wire  _T_1514; // @[util.scala 60:60:@3381.4]
  wire  _T_1515; // @[util.scala 60:60:@3382.4]
  wire  _T_1516; // @[util.scala 60:60:@3383.4]
  wire  _T_1517; // @[util.scala 60:60:@3384.4]
  wire  _T_1518; // @[util.scala 60:60:@3385.4]
  wire  _T_1519; // @[util.scala 60:60:@3386.4]
  wire  _T_1520; // @[util.scala 60:60:@3387.4]
  wire [255:0] _T_2299; // @[Mux.scala 19:72:@3839.4]
  wire [255:0] _T_2301; // @[Mux.scala 19:72:@3840.4]
  wire [255:0] _T_2308; // @[Mux.scala 19:72:@3847.4]
  wire [255:0] _T_2310; // @[Mux.scala 19:72:@3848.4]
  wire [255:0] _T_2317; // @[Mux.scala 19:72:@3855.4]
  wire [255:0] _T_2319; // @[Mux.scala 19:72:@3856.4]
  wire [255:0] _T_2326; // @[Mux.scala 19:72:@3863.4]
  wire [255:0] _T_2328; // @[Mux.scala 19:72:@3864.4]
  wire [255:0] _T_2335; // @[Mux.scala 19:72:@3871.4]
  wire [255:0] _T_2337; // @[Mux.scala 19:72:@3872.4]
  wire [255:0] _T_2344; // @[Mux.scala 19:72:@3879.4]
  wire [255:0] _T_2346; // @[Mux.scala 19:72:@3880.4]
  wire [255:0] _T_2353; // @[Mux.scala 19:72:@3887.4]
  wire [255:0] _T_2355; // @[Mux.scala 19:72:@3888.4]
  wire [255:0] _T_2362; // @[Mux.scala 19:72:@3895.4]
  wire [255:0] _T_2364; // @[Mux.scala 19:72:@3896.4]
  wire [255:0] _T_2365; // @[Mux.scala 19:72:@3897.4]
  wire [255:0] _T_2366; // @[Mux.scala 19:72:@3898.4]
  wire [255:0] _T_2367; // @[Mux.scala 19:72:@3899.4]
  wire [255:0] _T_2368; // @[Mux.scala 19:72:@3900.4]
  wire [255:0] _T_2369; // @[Mux.scala 19:72:@3901.4]
  wire [255:0] _T_2370; // @[Mux.scala 19:72:@3902.4]
  wire [255:0] _T_2371; // @[Mux.scala 19:72:@3903.4]
  wire [7:0] _T_2612; // @[Mux.scala 19:72:@4021.4]
  wire [7:0] _T_2614; // @[Mux.scala 19:72:@4022.4]
  wire [7:0] _T_2621; // @[Mux.scala 19:72:@4029.4]
  wire [7:0] _T_2623; // @[Mux.scala 19:72:@4030.4]
  wire [7:0] _T_2630; // @[Mux.scala 19:72:@4037.4]
  wire [7:0] _T_2632; // @[Mux.scala 19:72:@4038.4]
  wire [7:0] _T_2639; // @[Mux.scala 19:72:@4045.4]
  wire [7:0] _T_2641; // @[Mux.scala 19:72:@4046.4]
  wire [7:0] _T_2648; // @[Mux.scala 19:72:@4053.4]
  wire [7:0] _T_2650; // @[Mux.scala 19:72:@4054.4]
  wire [7:0] _T_2657; // @[Mux.scala 19:72:@4061.4]
  wire [7:0] _T_2659; // @[Mux.scala 19:72:@4062.4]
  wire [7:0] _T_2666; // @[Mux.scala 19:72:@4069.4]
  wire [7:0] _T_2668; // @[Mux.scala 19:72:@4070.4]
  wire [7:0] _T_2675; // @[Mux.scala 19:72:@4077.4]
  wire [7:0] _T_2677; // @[Mux.scala 19:72:@4078.4]
  wire [7:0] _T_2678; // @[Mux.scala 19:72:@4079.4]
  wire [7:0] _T_2679; // @[Mux.scala 19:72:@4080.4]
  wire [7:0] _T_2680; // @[Mux.scala 19:72:@4081.4]
  wire [7:0] _T_2681; // @[Mux.scala 19:72:@4082.4]
  wire [7:0] _T_2682; // @[Mux.scala 19:72:@4083.4]
  wire [7:0] _T_2683; // @[Mux.scala 19:72:@4084.4]
  wire [7:0] _T_2684; // @[Mux.scala 19:72:@4085.4]
  wire  _T_2761; // @[LoadQueue.scala 121:105:@4105.4]
  wire  _T_2763; // @[LoadQueue.scala 122:18:@4106.4]
  wire  _T_2765; // @[LoadQueue.scala 122:36:@4107.4]
  wire  _T_2766; // @[LoadQueue.scala 122:27:@4108.4]
  wire  _T_2768; // @[LoadQueue.scala 122:52:@4109.4]
  wire  _T_2770; // @[LoadQueue.scala 122:85:@4110.4]
  wire  _T_2772; // @[LoadQueue.scala 122:103:@4111.4]
  wire  _T_2773; // @[LoadQueue.scala 122:94:@4112.4]
  wire  _T_2775; // @[LoadQueue.scala 122:70:@4113.4]
  wire  _T_2776; // @[LoadQueue.scala 122:67:@4114.4]
  wire  validEntriesInStoreQ_0; // @[LoadQueue.scala 121:91:@4115.4]
  wire  _T_2780; // @[LoadQueue.scala 122:18:@4117.4]
  wire  _T_2782; // @[LoadQueue.scala 122:36:@4118.4]
  wire  _T_2783; // @[LoadQueue.scala 122:27:@4119.4]
  wire  _T_2787; // @[LoadQueue.scala 122:85:@4121.4]
  wire  _T_2789; // @[LoadQueue.scala 122:103:@4122.4]
  wire  _T_2790; // @[LoadQueue.scala 122:94:@4123.4]
  wire  _T_2792; // @[LoadQueue.scala 122:70:@4124.4]
  wire  _T_2793; // @[LoadQueue.scala 122:67:@4125.4]
  wire  validEntriesInStoreQ_1; // @[LoadQueue.scala 121:91:@4126.4]
  wire  _T_2797; // @[LoadQueue.scala 122:18:@4128.4]
  wire  _T_2799; // @[LoadQueue.scala 122:36:@4129.4]
  wire  _T_2800; // @[LoadQueue.scala 122:27:@4130.4]
  wire  _T_2804; // @[LoadQueue.scala 122:85:@4132.4]
  wire  _T_2806; // @[LoadQueue.scala 122:103:@4133.4]
  wire  _T_2807; // @[LoadQueue.scala 122:94:@4134.4]
  wire  _T_2809; // @[LoadQueue.scala 122:70:@4135.4]
  wire  _T_2810; // @[LoadQueue.scala 122:67:@4136.4]
  wire  validEntriesInStoreQ_2; // @[LoadQueue.scala 121:91:@4137.4]
  wire  _T_2814; // @[LoadQueue.scala 122:18:@4139.4]
  wire  _T_2816; // @[LoadQueue.scala 122:36:@4140.4]
  wire  _T_2817; // @[LoadQueue.scala 122:27:@4141.4]
  wire  _T_2821; // @[LoadQueue.scala 122:85:@4143.4]
  wire  _T_2823; // @[LoadQueue.scala 122:103:@4144.4]
  wire  _T_2824; // @[LoadQueue.scala 122:94:@4145.4]
  wire  _T_2826; // @[LoadQueue.scala 122:70:@4146.4]
  wire  _T_2827; // @[LoadQueue.scala 122:67:@4147.4]
  wire  validEntriesInStoreQ_3; // @[LoadQueue.scala 121:91:@4148.4]
  wire  _T_2831; // @[LoadQueue.scala 122:18:@4150.4]
  wire  _T_2833; // @[LoadQueue.scala 122:36:@4151.4]
  wire  _T_2834; // @[LoadQueue.scala 122:27:@4152.4]
  wire  _T_2838; // @[LoadQueue.scala 122:85:@4154.4]
  wire  _T_2840; // @[LoadQueue.scala 122:103:@4155.4]
  wire  _T_2841; // @[LoadQueue.scala 122:94:@4156.4]
  wire  _T_2843; // @[LoadQueue.scala 122:70:@4157.4]
  wire  _T_2844; // @[LoadQueue.scala 122:67:@4158.4]
  wire  validEntriesInStoreQ_4; // @[LoadQueue.scala 121:91:@4159.4]
  wire  _T_2848; // @[LoadQueue.scala 122:18:@4161.4]
  wire  _T_2850; // @[LoadQueue.scala 122:36:@4162.4]
  wire  _T_2851; // @[LoadQueue.scala 122:27:@4163.4]
  wire  _T_2855; // @[LoadQueue.scala 122:85:@4165.4]
  wire  _T_2857; // @[LoadQueue.scala 122:103:@4166.4]
  wire  _T_2858; // @[LoadQueue.scala 122:94:@4167.4]
  wire  _T_2860; // @[LoadQueue.scala 122:70:@4168.4]
  wire  _T_2861; // @[LoadQueue.scala 122:67:@4169.4]
  wire  validEntriesInStoreQ_5; // @[LoadQueue.scala 121:91:@4170.4]
  wire  _T_2865; // @[LoadQueue.scala 122:18:@4172.4]
  wire  _T_2867; // @[LoadQueue.scala 122:36:@4173.4]
  wire  _T_2868; // @[LoadQueue.scala 122:27:@4174.4]
  wire  _T_2872; // @[LoadQueue.scala 122:85:@4176.4]
  wire  _T_2874; // @[LoadQueue.scala 122:103:@4177.4]
  wire  _T_2875; // @[LoadQueue.scala 122:94:@4178.4]
  wire  _T_2877; // @[LoadQueue.scala 122:70:@4179.4]
  wire  _T_2878; // @[LoadQueue.scala 122:67:@4180.4]
  wire  validEntriesInStoreQ_6; // @[LoadQueue.scala 121:91:@4181.4]
  wire  validEntriesInStoreQ_7; // @[LoadQueue.scala 121:91:@4192.4]
  wire  storesToCheck_0_0; // @[LoadQueue.scala 131:10:@4211.4]
  wire  _T_3294; // @[LoadQueue.scala 131:81:@4214.4]
  wire  _T_3295; // @[LoadQueue.scala 131:72:@4215.4]
  wire  _T_3297; // @[LoadQueue.scala 132:33:@4216.4]
  wire  _T_3300; // @[LoadQueue.scala 132:41:@4218.4]
  wire  _T_3302; // @[LoadQueue.scala 132:9:@4219.4]
  wire  storesToCheck_0_1; // @[LoadQueue.scala 131:10:@4220.4]
  wire  _T_3308; // @[LoadQueue.scala 131:81:@4223.4]
  wire  _T_3309; // @[LoadQueue.scala 131:72:@4224.4]
  wire  _T_3311; // @[LoadQueue.scala 132:33:@4225.4]
  wire  _T_3314; // @[LoadQueue.scala 132:41:@4227.4]
  wire  _T_3316; // @[LoadQueue.scala 132:9:@4228.4]
  wire  storesToCheck_0_2; // @[LoadQueue.scala 131:10:@4229.4]
  wire  _T_3322; // @[LoadQueue.scala 131:81:@4232.4]
  wire  _T_3323; // @[LoadQueue.scala 131:72:@4233.4]
  wire  _T_3325; // @[LoadQueue.scala 132:33:@4234.4]
  wire  _T_3328; // @[LoadQueue.scala 132:41:@4236.4]
  wire  _T_3330; // @[LoadQueue.scala 132:9:@4237.4]
  wire  storesToCheck_0_3; // @[LoadQueue.scala 131:10:@4238.4]
  wire  _T_3336; // @[LoadQueue.scala 131:81:@4241.4]
  wire  _T_3337; // @[LoadQueue.scala 131:72:@4242.4]
  wire  _T_3339; // @[LoadQueue.scala 132:33:@4243.4]
  wire  _T_3342; // @[LoadQueue.scala 132:41:@4245.4]
  wire  _T_3344; // @[LoadQueue.scala 132:9:@4246.4]
  wire  storesToCheck_0_4; // @[LoadQueue.scala 131:10:@4247.4]
  wire  _T_3350; // @[LoadQueue.scala 131:81:@4250.4]
  wire  _T_3351; // @[LoadQueue.scala 131:72:@4251.4]
  wire  _T_3353; // @[LoadQueue.scala 132:33:@4252.4]
  wire  _T_3356; // @[LoadQueue.scala 132:41:@4254.4]
  wire  _T_3358; // @[LoadQueue.scala 132:9:@4255.4]
  wire  storesToCheck_0_5; // @[LoadQueue.scala 131:10:@4256.4]
  wire  _T_3364; // @[LoadQueue.scala 131:81:@4259.4]
  wire  _T_3365; // @[LoadQueue.scala 131:72:@4260.4]
  wire  _T_3367; // @[LoadQueue.scala 132:33:@4261.4]
  wire  _T_3370; // @[LoadQueue.scala 132:41:@4263.4]
  wire  _T_3372; // @[LoadQueue.scala 132:9:@4264.4]
  wire  storesToCheck_0_6; // @[LoadQueue.scala 131:10:@4265.4]
  wire  _T_3378; // @[LoadQueue.scala 131:81:@4268.4]
  wire  storesToCheck_0_7; // @[LoadQueue.scala 131:10:@4274.4]
  wire  storesToCheck_1_0; // @[LoadQueue.scala 131:10:@4300.4]
  wire  _T_3420; // @[LoadQueue.scala 131:81:@4303.4]
  wire  _T_3421; // @[LoadQueue.scala 131:72:@4304.4]
  wire  _T_3423; // @[LoadQueue.scala 132:33:@4305.4]
  wire  _T_3426; // @[LoadQueue.scala 132:41:@4307.4]
  wire  _T_3428; // @[LoadQueue.scala 132:9:@4308.4]
  wire  storesToCheck_1_1; // @[LoadQueue.scala 131:10:@4309.4]
  wire  _T_3434; // @[LoadQueue.scala 131:81:@4312.4]
  wire  _T_3435; // @[LoadQueue.scala 131:72:@4313.4]
  wire  _T_3437; // @[LoadQueue.scala 132:33:@4314.4]
  wire  _T_3440; // @[LoadQueue.scala 132:41:@4316.4]
  wire  _T_3442; // @[LoadQueue.scala 132:9:@4317.4]
  wire  storesToCheck_1_2; // @[LoadQueue.scala 131:10:@4318.4]
  wire  _T_3448; // @[LoadQueue.scala 131:81:@4321.4]
  wire  _T_3449; // @[LoadQueue.scala 131:72:@4322.4]
  wire  _T_3451; // @[LoadQueue.scala 132:33:@4323.4]
  wire  _T_3454; // @[LoadQueue.scala 132:41:@4325.4]
  wire  _T_3456; // @[LoadQueue.scala 132:9:@4326.4]
  wire  storesToCheck_1_3; // @[LoadQueue.scala 131:10:@4327.4]
  wire  _T_3462; // @[LoadQueue.scala 131:81:@4330.4]
  wire  _T_3463; // @[LoadQueue.scala 131:72:@4331.4]
  wire  _T_3465; // @[LoadQueue.scala 132:33:@4332.4]
  wire  _T_3468; // @[LoadQueue.scala 132:41:@4334.4]
  wire  _T_3470; // @[LoadQueue.scala 132:9:@4335.4]
  wire  storesToCheck_1_4; // @[LoadQueue.scala 131:10:@4336.4]
  wire  _T_3476; // @[LoadQueue.scala 131:81:@4339.4]
  wire  _T_3477; // @[LoadQueue.scala 131:72:@4340.4]
  wire  _T_3479; // @[LoadQueue.scala 132:33:@4341.4]
  wire  _T_3482; // @[LoadQueue.scala 132:41:@4343.4]
  wire  _T_3484; // @[LoadQueue.scala 132:9:@4344.4]
  wire  storesToCheck_1_5; // @[LoadQueue.scala 131:10:@4345.4]
  wire  _T_3490; // @[LoadQueue.scala 131:81:@4348.4]
  wire  _T_3491; // @[LoadQueue.scala 131:72:@4349.4]
  wire  _T_3493; // @[LoadQueue.scala 132:33:@4350.4]
  wire  _T_3496; // @[LoadQueue.scala 132:41:@4352.4]
  wire  _T_3498; // @[LoadQueue.scala 132:9:@4353.4]
  wire  storesToCheck_1_6; // @[LoadQueue.scala 131:10:@4354.4]
  wire  _T_3504; // @[LoadQueue.scala 131:81:@4357.4]
  wire  storesToCheck_1_7; // @[LoadQueue.scala 131:10:@4363.4]
  wire  storesToCheck_2_0; // @[LoadQueue.scala 131:10:@4389.4]
  wire  _T_3546; // @[LoadQueue.scala 131:81:@4392.4]
  wire  _T_3547; // @[LoadQueue.scala 131:72:@4393.4]
  wire  _T_3549; // @[LoadQueue.scala 132:33:@4394.4]
  wire  _T_3552; // @[LoadQueue.scala 132:41:@4396.4]
  wire  _T_3554; // @[LoadQueue.scala 132:9:@4397.4]
  wire  storesToCheck_2_1; // @[LoadQueue.scala 131:10:@4398.4]
  wire  _T_3560; // @[LoadQueue.scala 131:81:@4401.4]
  wire  _T_3561; // @[LoadQueue.scala 131:72:@4402.4]
  wire  _T_3563; // @[LoadQueue.scala 132:33:@4403.4]
  wire  _T_3566; // @[LoadQueue.scala 132:41:@4405.4]
  wire  _T_3568; // @[LoadQueue.scala 132:9:@4406.4]
  wire  storesToCheck_2_2; // @[LoadQueue.scala 131:10:@4407.4]
  wire  _T_3574; // @[LoadQueue.scala 131:81:@4410.4]
  wire  _T_3575; // @[LoadQueue.scala 131:72:@4411.4]
  wire  _T_3577; // @[LoadQueue.scala 132:33:@4412.4]
  wire  _T_3580; // @[LoadQueue.scala 132:41:@4414.4]
  wire  _T_3582; // @[LoadQueue.scala 132:9:@4415.4]
  wire  storesToCheck_2_3; // @[LoadQueue.scala 131:10:@4416.4]
  wire  _T_3588; // @[LoadQueue.scala 131:81:@4419.4]
  wire  _T_3589; // @[LoadQueue.scala 131:72:@4420.4]
  wire  _T_3591; // @[LoadQueue.scala 132:33:@4421.4]
  wire  _T_3594; // @[LoadQueue.scala 132:41:@4423.4]
  wire  _T_3596; // @[LoadQueue.scala 132:9:@4424.4]
  wire  storesToCheck_2_4; // @[LoadQueue.scala 131:10:@4425.4]
  wire  _T_3602; // @[LoadQueue.scala 131:81:@4428.4]
  wire  _T_3603; // @[LoadQueue.scala 131:72:@4429.4]
  wire  _T_3605; // @[LoadQueue.scala 132:33:@4430.4]
  wire  _T_3608; // @[LoadQueue.scala 132:41:@4432.4]
  wire  _T_3610; // @[LoadQueue.scala 132:9:@4433.4]
  wire  storesToCheck_2_5; // @[LoadQueue.scala 131:10:@4434.4]
  wire  _T_3616; // @[LoadQueue.scala 131:81:@4437.4]
  wire  _T_3617; // @[LoadQueue.scala 131:72:@4438.4]
  wire  _T_3619; // @[LoadQueue.scala 132:33:@4439.4]
  wire  _T_3622; // @[LoadQueue.scala 132:41:@4441.4]
  wire  _T_3624; // @[LoadQueue.scala 132:9:@4442.4]
  wire  storesToCheck_2_6; // @[LoadQueue.scala 131:10:@4443.4]
  wire  _T_3630; // @[LoadQueue.scala 131:81:@4446.4]
  wire  storesToCheck_2_7; // @[LoadQueue.scala 131:10:@4452.4]
  wire  storesToCheck_3_0; // @[LoadQueue.scala 131:10:@4478.4]
  wire  _T_3672; // @[LoadQueue.scala 131:81:@4481.4]
  wire  _T_3673; // @[LoadQueue.scala 131:72:@4482.4]
  wire  _T_3675; // @[LoadQueue.scala 132:33:@4483.4]
  wire  _T_3678; // @[LoadQueue.scala 132:41:@4485.4]
  wire  _T_3680; // @[LoadQueue.scala 132:9:@4486.4]
  wire  storesToCheck_3_1; // @[LoadQueue.scala 131:10:@4487.4]
  wire  _T_3686; // @[LoadQueue.scala 131:81:@4490.4]
  wire  _T_3687; // @[LoadQueue.scala 131:72:@4491.4]
  wire  _T_3689; // @[LoadQueue.scala 132:33:@4492.4]
  wire  _T_3692; // @[LoadQueue.scala 132:41:@4494.4]
  wire  _T_3694; // @[LoadQueue.scala 132:9:@4495.4]
  wire  storesToCheck_3_2; // @[LoadQueue.scala 131:10:@4496.4]
  wire  _T_3700; // @[LoadQueue.scala 131:81:@4499.4]
  wire  _T_3701; // @[LoadQueue.scala 131:72:@4500.4]
  wire  _T_3703; // @[LoadQueue.scala 132:33:@4501.4]
  wire  _T_3706; // @[LoadQueue.scala 132:41:@4503.4]
  wire  _T_3708; // @[LoadQueue.scala 132:9:@4504.4]
  wire  storesToCheck_3_3; // @[LoadQueue.scala 131:10:@4505.4]
  wire  _T_3714; // @[LoadQueue.scala 131:81:@4508.4]
  wire  _T_3715; // @[LoadQueue.scala 131:72:@4509.4]
  wire  _T_3717; // @[LoadQueue.scala 132:33:@4510.4]
  wire  _T_3720; // @[LoadQueue.scala 132:41:@4512.4]
  wire  _T_3722; // @[LoadQueue.scala 132:9:@4513.4]
  wire  storesToCheck_3_4; // @[LoadQueue.scala 131:10:@4514.4]
  wire  _T_3728; // @[LoadQueue.scala 131:81:@4517.4]
  wire  _T_3729; // @[LoadQueue.scala 131:72:@4518.4]
  wire  _T_3731; // @[LoadQueue.scala 132:33:@4519.4]
  wire  _T_3734; // @[LoadQueue.scala 132:41:@4521.4]
  wire  _T_3736; // @[LoadQueue.scala 132:9:@4522.4]
  wire  storesToCheck_3_5; // @[LoadQueue.scala 131:10:@4523.4]
  wire  _T_3742; // @[LoadQueue.scala 131:81:@4526.4]
  wire  _T_3743; // @[LoadQueue.scala 131:72:@4527.4]
  wire  _T_3745; // @[LoadQueue.scala 132:33:@4528.4]
  wire  _T_3748; // @[LoadQueue.scala 132:41:@4530.4]
  wire  _T_3750; // @[LoadQueue.scala 132:9:@4531.4]
  wire  storesToCheck_3_6; // @[LoadQueue.scala 131:10:@4532.4]
  wire  _T_3756; // @[LoadQueue.scala 131:81:@4535.4]
  wire  storesToCheck_3_7; // @[LoadQueue.scala 131:10:@4541.4]
  wire  storesToCheck_4_0; // @[LoadQueue.scala 131:10:@4567.4]
  wire  _T_3798; // @[LoadQueue.scala 131:81:@4570.4]
  wire  _T_3799; // @[LoadQueue.scala 131:72:@4571.4]
  wire  _T_3801; // @[LoadQueue.scala 132:33:@4572.4]
  wire  _T_3804; // @[LoadQueue.scala 132:41:@4574.4]
  wire  _T_3806; // @[LoadQueue.scala 132:9:@4575.4]
  wire  storesToCheck_4_1; // @[LoadQueue.scala 131:10:@4576.4]
  wire  _T_3812; // @[LoadQueue.scala 131:81:@4579.4]
  wire  _T_3813; // @[LoadQueue.scala 131:72:@4580.4]
  wire  _T_3815; // @[LoadQueue.scala 132:33:@4581.4]
  wire  _T_3818; // @[LoadQueue.scala 132:41:@4583.4]
  wire  _T_3820; // @[LoadQueue.scala 132:9:@4584.4]
  wire  storesToCheck_4_2; // @[LoadQueue.scala 131:10:@4585.4]
  wire  _T_3826; // @[LoadQueue.scala 131:81:@4588.4]
  wire  _T_3827; // @[LoadQueue.scala 131:72:@4589.4]
  wire  _T_3829; // @[LoadQueue.scala 132:33:@4590.4]
  wire  _T_3832; // @[LoadQueue.scala 132:41:@4592.4]
  wire  _T_3834; // @[LoadQueue.scala 132:9:@4593.4]
  wire  storesToCheck_4_3; // @[LoadQueue.scala 131:10:@4594.4]
  wire  _T_3840; // @[LoadQueue.scala 131:81:@4597.4]
  wire  _T_3841; // @[LoadQueue.scala 131:72:@4598.4]
  wire  _T_3843; // @[LoadQueue.scala 132:33:@4599.4]
  wire  _T_3846; // @[LoadQueue.scala 132:41:@4601.4]
  wire  _T_3848; // @[LoadQueue.scala 132:9:@4602.4]
  wire  storesToCheck_4_4; // @[LoadQueue.scala 131:10:@4603.4]
  wire  _T_3854; // @[LoadQueue.scala 131:81:@4606.4]
  wire  _T_3855; // @[LoadQueue.scala 131:72:@4607.4]
  wire  _T_3857; // @[LoadQueue.scala 132:33:@4608.4]
  wire  _T_3860; // @[LoadQueue.scala 132:41:@4610.4]
  wire  _T_3862; // @[LoadQueue.scala 132:9:@4611.4]
  wire  storesToCheck_4_5; // @[LoadQueue.scala 131:10:@4612.4]
  wire  _T_3868; // @[LoadQueue.scala 131:81:@4615.4]
  wire  _T_3869; // @[LoadQueue.scala 131:72:@4616.4]
  wire  _T_3871; // @[LoadQueue.scala 132:33:@4617.4]
  wire  _T_3874; // @[LoadQueue.scala 132:41:@4619.4]
  wire  _T_3876; // @[LoadQueue.scala 132:9:@4620.4]
  wire  storesToCheck_4_6; // @[LoadQueue.scala 131:10:@4621.4]
  wire  _T_3882; // @[LoadQueue.scala 131:81:@4624.4]
  wire  storesToCheck_4_7; // @[LoadQueue.scala 131:10:@4630.4]
  wire  storesToCheck_5_0; // @[LoadQueue.scala 131:10:@4656.4]
  wire  _T_3924; // @[LoadQueue.scala 131:81:@4659.4]
  wire  _T_3925; // @[LoadQueue.scala 131:72:@4660.4]
  wire  _T_3927; // @[LoadQueue.scala 132:33:@4661.4]
  wire  _T_3930; // @[LoadQueue.scala 132:41:@4663.4]
  wire  _T_3932; // @[LoadQueue.scala 132:9:@4664.4]
  wire  storesToCheck_5_1; // @[LoadQueue.scala 131:10:@4665.4]
  wire  _T_3938; // @[LoadQueue.scala 131:81:@4668.4]
  wire  _T_3939; // @[LoadQueue.scala 131:72:@4669.4]
  wire  _T_3941; // @[LoadQueue.scala 132:33:@4670.4]
  wire  _T_3944; // @[LoadQueue.scala 132:41:@4672.4]
  wire  _T_3946; // @[LoadQueue.scala 132:9:@4673.4]
  wire  storesToCheck_5_2; // @[LoadQueue.scala 131:10:@4674.4]
  wire  _T_3952; // @[LoadQueue.scala 131:81:@4677.4]
  wire  _T_3953; // @[LoadQueue.scala 131:72:@4678.4]
  wire  _T_3955; // @[LoadQueue.scala 132:33:@4679.4]
  wire  _T_3958; // @[LoadQueue.scala 132:41:@4681.4]
  wire  _T_3960; // @[LoadQueue.scala 132:9:@4682.4]
  wire  storesToCheck_5_3; // @[LoadQueue.scala 131:10:@4683.4]
  wire  _T_3966; // @[LoadQueue.scala 131:81:@4686.4]
  wire  _T_3967; // @[LoadQueue.scala 131:72:@4687.4]
  wire  _T_3969; // @[LoadQueue.scala 132:33:@4688.4]
  wire  _T_3972; // @[LoadQueue.scala 132:41:@4690.4]
  wire  _T_3974; // @[LoadQueue.scala 132:9:@4691.4]
  wire  storesToCheck_5_4; // @[LoadQueue.scala 131:10:@4692.4]
  wire  _T_3980; // @[LoadQueue.scala 131:81:@4695.4]
  wire  _T_3981; // @[LoadQueue.scala 131:72:@4696.4]
  wire  _T_3983; // @[LoadQueue.scala 132:33:@4697.4]
  wire  _T_3986; // @[LoadQueue.scala 132:41:@4699.4]
  wire  _T_3988; // @[LoadQueue.scala 132:9:@4700.4]
  wire  storesToCheck_5_5; // @[LoadQueue.scala 131:10:@4701.4]
  wire  _T_3994; // @[LoadQueue.scala 131:81:@4704.4]
  wire  _T_3995; // @[LoadQueue.scala 131:72:@4705.4]
  wire  _T_3997; // @[LoadQueue.scala 132:33:@4706.4]
  wire  _T_4000; // @[LoadQueue.scala 132:41:@4708.4]
  wire  _T_4002; // @[LoadQueue.scala 132:9:@4709.4]
  wire  storesToCheck_5_6; // @[LoadQueue.scala 131:10:@4710.4]
  wire  _T_4008; // @[LoadQueue.scala 131:81:@4713.4]
  wire  storesToCheck_5_7; // @[LoadQueue.scala 131:10:@4719.4]
  wire  storesToCheck_6_0; // @[LoadQueue.scala 131:10:@4745.4]
  wire  _T_4050; // @[LoadQueue.scala 131:81:@4748.4]
  wire  _T_4051; // @[LoadQueue.scala 131:72:@4749.4]
  wire  _T_4053; // @[LoadQueue.scala 132:33:@4750.4]
  wire  _T_4056; // @[LoadQueue.scala 132:41:@4752.4]
  wire  _T_4058; // @[LoadQueue.scala 132:9:@4753.4]
  wire  storesToCheck_6_1; // @[LoadQueue.scala 131:10:@4754.4]
  wire  _T_4064; // @[LoadQueue.scala 131:81:@4757.4]
  wire  _T_4065; // @[LoadQueue.scala 131:72:@4758.4]
  wire  _T_4067; // @[LoadQueue.scala 132:33:@4759.4]
  wire  _T_4070; // @[LoadQueue.scala 132:41:@4761.4]
  wire  _T_4072; // @[LoadQueue.scala 132:9:@4762.4]
  wire  storesToCheck_6_2; // @[LoadQueue.scala 131:10:@4763.4]
  wire  _T_4078; // @[LoadQueue.scala 131:81:@4766.4]
  wire  _T_4079; // @[LoadQueue.scala 131:72:@4767.4]
  wire  _T_4081; // @[LoadQueue.scala 132:33:@4768.4]
  wire  _T_4084; // @[LoadQueue.scala 132:41:@4770.4]
  wire  _T_4086; // @[LoadQueue.scala 132:9:@4771.4]
  wire  storesToCheck_6_3; // @[LoadQueue.scala 131:10:@4772.4]
  wire  _T_4092; // @[LoadQueue.scala 131:81:@4775.4]
  wire  _T_4093; // @[LoadQueue.scala 131:72:@4776.4]
  wire  _T_4095; // @[LoadQueue.scala 132:33:@4777.4]
  wire  _T_4098; // @[LoadQueue.scala 132:41:@4779.4]
  wire  _T_4100; // @[LoadQueue.scala 132:9:@4780.4]
  wire  storesToCheck_6_4; // @[LoadQueue.scala 131:10:@4781.4]
  wire  _T_4106; // @[LoadQueue.scala 131:81:@4784.4]
  wire  _T_4107; // @[LoadQueue.scala 131:72:@4785.4]
  wire  _T_4109; // @[LoadQueue.scala 132:33:@4786.4]
  wire  _T_4112; // @[LoadQueue.scala 132:41:@4788.4]
  wire  _T_4114; // @[LoadQueue.scala 132:9:@4789.4]
  wire  storesToCheck_6_5; // @[LoadQueue.scala 131:10:@4790.4]
  wire  _T_4120; // @[LoadQueue.scala 131:81:@4793.4]
  wire  _T_4121; // @[LoadQueue.scala 131:72:@4794.4]
  wire  _T_4123; // @[LoadQueue.scala 132:33:@4795.4]
  wire  _T_4126; // @[LoadQueue.scala 132:41:@4797.4]
  wire  _T_4128; // @[LoadQueue.scala 132:9:@4798.4]
  wire  storesToCheck_6_6; // @[LoadQueue.scala 131:10:@4799.4]
  wire  _T_4134; // @[LoadQueue.scala 131:81:@4802.4]
  wire  storesToCheck_6_7; // @[LoadQueue.scala 131:10:@4808.4]
  wire  storesToCheck_7_0; // @[LoadQueue.scala 131:10:@4834.4]
  wire  _T_4176; // @[LoadQueue.scala 131:81:@4837.4]
  wire  _T_4177; // @[LoadQueue.scala 131:72:@4838.4]
  wire  _T_4179; // @[LoadQueue.scala 132:33:@4839.4]
  wire  _T_4182; // @[LoadQueue.scala 132:41:@4841.4]
  wire  _T_4184; // @[LoadQueue.scala 132:9:@4842.4]
  wire  storesToCheck_7_1; // @[LoadQueue.scala 131:10:@4843.4]
  wire  _T_4190; // @[LoadQueue.scala 131:81:@4846.4]
  wire  _T_4191; // @[LoadQueue.scala 131:72:@4847.4]
  wire  _T_4193; // @[LoadQueue.scala 132:33:@4848.4]
  wire  _T_4196; // @[LoadQueue.scala 132:41:@4850.4]
  wire  _T_4198; // @[LoadQueue.scala 132:9:@4851.4]
  wire  storesToCheck_7_2; // @[LoadQueue.scala 131:10:@4852.4]
  wire  _T_4204; // @[LoadQueue.scala 131:81:@4855.4]
  wire  _T_4205; // @[LoadQueue.scala 131:72:@4856.4]
  wire  _T_4207; // @[LoadQueue.scala 132:33:@4857.4]
  wire  _T_4210; // @[LoadQueue.scala 132:41:@4859.4]
  wire  _T_4212; // @[LoadQueue.scala 132:9:@4860.4]
  wire  storesToCheck_7_3; // @[LoadQueue.scala 131:10:@4861.4]
  wire  _T_4218; // @[LoadQueue.scala 131:81:@4864.4]
  wire  _T_4219; // @[LoadQueue.scala 131:72:@4865.4]
  wire  _T_4221; // @[LoadQueue.scala 132:33:@4866.4]
  wire  _T_4224; // @[LoadQueue.scala 132:41:@4868.4]
  wire  _T_4226; // @[LoadQueue.scala 132:9:@4869.4]
  wire  storesToCheck_7_4; // @[LoadQueue.scala 131:10:@4870.4]
  wire  _T_4232; // @[LoadQueue.scala 131:81:@4873.4]
  wire  _T_4233; // @[LoadQueue.scala 131:72:@4874.4]
  wire  _T_4235; // @[LoadQueue.scala 132:33:@4875.4]
  wire  _T_4238; // @[LoadQueue.scala 132:41:@4877.4]
  wire  _T_4240; // @[LoadQueue.scala 132:9:@4878.4]
  wire  storesToCheck_7_5; // @[LoadQueue.scala 131:10:@4879.4]
  wire  _T_4246; // @[LoadQueue.scala 131:81:@4882.4]
  wire  _T_4247; // @[LoadQueue.scala 131:72:@4883.4]
  wire  _T_4249; // @[LoadQueue.scala 132:33:@4884.4]
  wire  _T_4252; // @[LoadQueue.scala 132:41:@4886.4]
  wire  _T_4254; // @[LoadQueue.scala 132:9:@4887.4]
  wire  storesToCheck_7_6; // @[LoadQueue.scala 131:10:@4888.4]
  wire  _T_4260; // @[LoadQueue.scala 131:81:@4891.4]
  wire  storesToCheck_7_7; // @[LoadQueue.scala 131:10:@4897.4]
  wire  _T_4650; // @[LoadQueue.scala 141:18:@4916.4]
  wire  entriesToCheck_0_0; // @[LoadQueue.scala 141:26:@4917.4]
  wire  _T_4652; // @[LoadQueue.scala 141:18:@4918.4]
  wire  entriesToCheck_0_1; // @[LoadQueue.scala 141:26:@4919.4]
  wire  _T_4654; // @[LoadQueue.scala 141:18:@4920.4]
  wire  entriesToCheck_0_2; // @[LoadQueue.scala 141:26:@4921.4]
  wire  _T_4656; // @[LoadQueue.scala 141:18:@4922.4]
  wire  entriesToCheck_0_3; // @[LoadQueue.scala 141:26:@4923.4]
  wire  _T_4658; // @[LoadQueue.scala 141:18:@4924.4]
  wire  entriesToCheck_0_4; // @[LoadQueue.scala 141:26:@4925.4]
  wire  _T_4660; // @[LoadQueue.scala 141:18:@4926.4]
  wire  entriesToCheck_0_5; // @[LoadQueue.scala 141:26:@4927.4]
  wire  _T_4662; // @[LoadQueue.scala 141:18:@4928.4]
  wire  entriesToCheck_0_6; // @[LoadQueue.scala 141:26:@4929.4]
  wire  _T_4664; // @[LoadQueue.scala 141:18:@4930.4]
  wire  entriesToCheck_0_7; // @[LoadQueue.scala 141:26:@4931.4]
  wire  _T_4666; // @[LoadQueue.scala 141:18:@4940.4]
  wire  entriesToCheck_1_0; // @[LoadQueue.scala 141:26:@4941.4]
  wire  _T_4668; // @[LoadQueue.scala 141:18:@4942.4]
  wire  entriesToCheck_1_1; // @[LoadQueue.scala 141:26:@4943.4]
  wire  _T_4670; // @[LoadQueue.scala 141:18:@4944.4]
  wire  entriesToCheck_1_2; // @[LoadQueue.scala 141:26:@4945.4]
  wire  _T_4672; // @[LoadQueue.scala 141:18:@4946.4]
  wire  entriesToCheck_1_3; // @[LoadQueue.scala 141:26:@4947.4]
  wire  _T_4674; // @[LoadQueue.scala 141:18:@4948.4]
  wire  entriesToCheck_1_4; // @[LoadQueue.scala 141:26:@4949.4]
  wire  _T_4676; // @[LoadQueue.scala 141:18:@4950.4]
  wire  entriesToCheck_1_5; // @[LoadQueue.scala 141:26:@4951.4]
  wire  _T_4678; // @[LoadQueue.scala 141:18:@4952.4]
  wire  entriesToCheck_1_6; // @[LoadQueue.scala 141:26:@4953.4]
  wire  _T_4680; // @[LoadQueue.scala 141:18:@4954.4]
  wire  entriesToCheck_1_7; // @[LoadQueue.scala 141:26:@4955.4]
  wire  _T_4682; // @[LoadQueue.scala 141:18:@4964.4]
  wire  entriesToCheck_2_0; // @[LoadQueue.scala 141:26:@4965.4]
  wire  _T_4684; // @[LoadQueue.scala 141:18:@4966.4]
  wire  entriesToCheck_2_1; // @[LoadQueue.scala 141:26:@4967.4]
  wire  _T_4686; // @[LoadQueue.scala 141:18:@4968.4]
  wire  entriesToCheck_2_2; // @[LoadQueue.scala 141:26:@4969.4]
  wire  _T_4688; // @[LoadQueue.scala 141:18:@4970.4]
  wire  entriesToCheck_2_3; // @[LoadQueue.scala 141:26:@4971.4]
  wire  _T_4690; // @[LoadQueue.scala 141:18:@4972.4]
  wire  entriesToCheck_2_4; // @[LoadQueue.scala 141:26:@4973.4]
  wire  _T_4692; // @[LoadQueue.scala 141:18:@4974.4]
  wire  entriesToCheck_2_5; // @[LoadQueue.scala 141:26:@4975.4]
  wire  _T_4694; // @[LoadQueue.scala 141:18:@4976.4]
  wire  entriesToCheck_2_6; // @[LoadQueue.scala 141:26:@4977.4]
  wire  _T_4696; // @[LoadQueue.scala 141:18:@4978.4]
  wire  entriesToCheck_2_7; // @[LoadQueue.scala 141:26:@4979.4]
  wire  _T_4698; // @[LoadQueue.scala 141:18:@4988.4]
  wire  entriesToCheck_3_0; // @[LoadQueue.scala 141:26:@4989.4]
  wire  _T_4700; // @[LoadQueue.scala 141:18:@4990.4]
  wire  entriesToCheck_3_1; // @[LoadQueue.scala 141:26:@4991.4]
  wire  _T_4702; // @[LoadQueue.scala 141:18:@4992.4]
  wire  entriesToCheck_3_2; // @[LoadQueue.scala 141:26:@4993.4]
  wire  _T_4704; // @[LoadQueue.scala 141:18:@4994.4]
  wire  entriesToCheck_3_3; // @[LoadQueue.scala 141:26:@4995.4]
  wire  _T_4706; // @[LoadQueue.scala 141:18:@4996.4]
  wire  entriesToCheck_3_4; // @[LoadQueue.scala 141:26:@4997.4]
  wire  _T_4708; // @[LoadQueue.scala 141:18:@4998.4]
  wire  entriesToCheck_3_5; // @[LoadQueue.scala 141:26:@4999.4]
  wire  _T_4710; // @[LoadQueue.scala 141:18:@5000.4]
  wire  entriesToCheck_3_6; // @[LoadQueue.scala 141:26:@5001.4]
  wire  _T_4712; // @[LoadQueue.scala 141:18:@5002.4]
  wire  entriesToCheck_3_7; // @[LoadQueue.scala 141:26:@5003.4]
  wire  _T_4714; // @[LoadQueue.scala 141:18:@5012.4]
  wire  entriesToCheck_4_0; // @[LoadQueue.scala 141:26:@5013.4]
  wire  _T_4716; // @[LoadQueue.scala 141:18:@5014.4]
  wire  entriesToCheck_4_1; // @[LoadQueue.scala 141:26:@5015.4]
  wire  _T_4718; // @[LoadQueue.scala 141:18:@5016.4]
  wire  entriesToCheck_4_2; // @[LoadQueue.scala 141:26:@5017.4]
  wire  _T_4720; // @[LoadQueue.scala 141:18:@5018.4]
  wire  entriesToCheck_4_3; // @[LoadQueue.scala 141:26:@5019.4]
  wire  _T_4722; // @[LoadQueue.scala 141:18:@5020.4]
  wire  entriesToCheck_4_4; // @[LoadQueue.scala 141:26:@5021.4]
  wire  _T_4724; // @[LoadQueue.scala 141:18:@5022.4]
  wire  entriesToCheck_4_5; // @[LoadQueue.scala 141:26:@5023.4]
  wire  _T_4726; // @[LoadQueue.scala 141:18:@5024.4]
  wire  entriesToCheck_4_6; // @[LoadQueue.scala 141:26:@5025.4]
  wire  _T_4728; // @[LoadQueue.scala 141:18:@5026.4]
  wire  entriesToCheck_4_7; // @[LoadQueue.scala 141:26:@5027.4]
  wire  _T_4730; // @[LoadQueue.scala 141:18:@5036.4]
  wire  entriesToCheck_5_0; // @[LoadQueue.scala 141:26:@5037.4]
  wire  _T_4732; // @[LoadQueue.scala 141:18:@5038.4]
  wire  entriesToCheck_5_1; // @[LoadQueue.scala 141:26:@5039.4]
  wire  _T_4734; // @[LoadQueue.scala 141:18:@5040.4]
  wire  entriesToCheck_5_2; // @[LoadQueue.scala 141:26:@5041.4]
  wire  _T_4736; // @[LoadQueue.scala 141:18:@5042.4]
  wire  entriesToCheck_5_3; // @[LoadQueue.scala 141:26:@5043.4]
  wire  _T_4738; // @[LoadQueue.scala 141:18:@5044.4]
  wire  entriesToCheck_5_4; // @[LoadQueue.scala 141:26:@5045.4]
  wire  _T_4740; // @[LoadQueue.scala 141:18:@5046.4]
  wire  entriesToCheck_5_5; // @[LoadQueue.scala 141:26:@5047.4]
  wire  _T_4742; // @[LoadQueue.scala 141:18:@5048.4]
  wire  entriesToCheck_5_6; // @[LoadQueue.scala 141:26:@5049.4]
  wire  _T_4744; // @[LoadQueue.scala 141:18:@5050.4]
  wire  entriesToCheck_5_7; // @[LoadQueue.scala 141:26:@5051.4]
  wire  _T_4746; // @[LoadQueue.scala 141:18:@5060.4]
  wire  entriesToCheck_6_0; // @[LoadQueue.scala 141:26:@5061.4]
  wire  _T_4748; // @[LoadQueue.scala 141:18:@5062.4]
  wire  entriesToCheck_6_1; // @[LoadQueue.scala 141:26:@5063.4]
  wire  _T_4750; // @[LoadQueue.scala 141:18:@5064.4]
  wire  entriesToCheck_6_2; // @[LoadQueue.scala 141:26:@5065.4]
  wire  _T_4752; // @[LoadQueue.scala 141:18:@5066.4]
  wire  entriesToCheck_6_3; // @[LoadQueue.scala 141:26:@5067.4]
  wire  _T_4754; // @[LoadQueue.scala 141:18:@5068.4]
  wire  entriesToCheck_6_4; // @[LoadQueue.scala 141:26:@5069.4]
  wire  _T_4756; // @[LoadQueue.scala 141:18:@5070.4]
  wire  entriesToCheck_6_5; // @[LoadQueue.scala 141:26:@5071.4]
  wire  _T_4758; // @[LoadQueue.scala 141:18:@5072.4]
  wire  entriesToCheck_6_6; // @[LoadQueue.scala 141:26:@5073.4]
  wire  _T_4760; // @[LoadQueue.scala 141:18:@5074.4]
  wire  entriesToCheck_6_7; // @[LoadQueue.scala 141:26:@5075.4]
  wire  _T_4762; // @[LoadQueue.scala 141:18:@5084.4]
  wire  entriesToCheck_7_0; // @[LoadQueue.scala 141:26:@5085.4]
  wire  _T_4764; // @[LoadQueue.scala 141:18:@5086.4]
  wire  entriesToCheck_7_1; // @[LoadQueue.scala 141:26:@5087.4]
  wire  _T_4766; // @[LoadQueue.scala 141:18:@5088.4]
  wire  entriesToCheck_7_2; // @[LoadQueue.scala 141:26:@5089.4]
  wire  _T_4768; // @[LoadQueue.scala 141:18:@5090.4]
  wire  entriesToCheck_7_3; // @[LoadQueue.scala 141:26:@5091.4]
  wire  _T_4770; // @[LoadQueue.scala 141:18:@5092.4]
  wire  entriesToCheck_7_4; // @[LoadQueue.scala 141:26:@5093.4]
  wire  _T_4772; // @[LoadQueue.scala 141:18:@5094.4]
  wire  entriesToCheck_7_5; // @[LoadQueue.scala 141:26:@5095.4]
  wire  _T_4774; // @[LoadQueue.scala 141:18:@5096.4]
  wire  entriesToCheck_7_6; // @[LoadQueue.scala 141:26:@5097.4]
  wire  _T_4776; // @[LoadQueue.scala 141:18:@5098.4]
  wire  entriesToCheck_7_7; // @[LoadQueue.scala 141:26:@5099.4]
  wire  _T_5144; // @[LoadQueue.scala 151:92:@5109.4]
  wire  _T_5145; // @[LoadQueue.scala 152:41:@5110.4]
  wire  _T_5146; // @[LoadQueue.scala 153:30:@5111.4]
  wire  conflict_0_0; // @[LoadQueue.scala 152:68:@5112.4]
  wire  _T_5148; // @[LoadQueue.scala 151:92:@5114.4]
  wire  _T_5149; // @[LoadQueue.scala 152:41:@5115.4]
  wire  _T_5150; // @[LoadQueue.scala 153:30:@5116.4]
  wire  conflict_0_1; // @[LoadQueue.scala 152:68:@5117.4]
  wire  _T_5152; // @[LoadQueue.scala 151:92:@5119.4]
  wire  _T_5153; // @[LoadQueue.scala 152:41:@5120.4]
  wire  _T_5154; // @[LoadQueue.scala 153:30:@5121.4]
  wire  conflict_0_2; // @[LoadQueue.scala 152:68:@5122.4]
  wire  _T_5156; // @[LoadQueue.scala 151:92:@5124.4]
  wire  _T_5157; // @[LoadQueue.scala 152:41:@5125.4]
  wire  _T_5158; // @[LoadQueue.scala 153:30:@5126.4]
  wire  conflict_0_3; // @[LoadQueue.scala 152:68:@5127.4]
  wire  _T_5160; // @[LoadQueue.scala 151:92:@5129.4]
  wire  _T_5161; // @[LoadQueue.scala 152:41:@5130.4]
  wire  _T_5162; // @[LoadQueue.scala 153:30:@5131.4]
  wire  conflict_0_4; // @[LoadQueue.scala 152:68:@5132.4]
  wire  _T_5164; // @[LoadQueue.scala 151:92:@5134.4]
  wire  _T_5165; // @[LoadQueue.scala 152:41:@5135.4]
  wire  _T_5166; // @[LoadQueue.scala 153:30:@5136.4]
  wire  conflict_0_5; // @[LoadQueue.scala 152:68:@5137.4]
  wire  _T_5168; // @[LoadQueue.scala 151:92:@5139.4]
  wire  _T_5169; // @[LoadQueue.scala 152:41:@5140.4]
  wire  _T_5170; // @[LoadQueue.scala 153:30:@5141.4]
  wire  conflict_0_6; // @[LoadQueue.scala 152:68:@5142.4]
  wire  _T_5172; // @[LoadQueue.scala 151:92:@5144.4]
  wire  _T_5173; // @[LoadQueue.scala 152:41:@5145.4]
  wire  _T_5174; // @[LoadQueue.scala 153:30:@5146.4]
  wire  conflict_0_7; // @[LoadQueue.scala 152:68:@5147.4]
  wire  _T_5176; // @[LoadQueue.scala 151:92:@5149.4]
  wire  _T_5177; // @[LoadQueue.scala 152:41:@5150.4]
  wire  _T_5178; // @[LoadQueue.scala 153:30:@5151.4]
  wire  conflict_1_0; // @[LoadQueue.scala 152:68:@5152.4]
  wire  _T_5180; // @[LoadQueue.scala 151:92:@5154.4]
  wire  _T_5181; // @[LoadQueue.scala 152:41:@5155.4]
  wire  _T_5182; // @[LoadQueue.scala 153:30:@5156.4]
  wire  conflict_1_1; // @[LoadQueue.scala 152:68:@5157.4]
  wire  _T_5184; // @[LoadQueue.scala 151:92:@5159.4]
  wire  _T_5185; // @[LoadQueue.scala 152:41:@5160.4]
  wire  _T_5186; // @[LoadQueue.scala 153:30:@5161.4]
  wire  conflict_1_2; // @[LoadQueue.scala 152:68:@5162.4]
  wire  _T_5188; // @[LoadQueue.scala 151:92:@5164.4]
  wire  _T_5189; // @[LoadQueue.scala 152:41:@5165.4]
  wire  _T_5190; // @[LoadQueue.scala 153:30:@5166.4]
  wire  conflict_1_3; // @[LoadQueue.scala 152:68:@5167.4]
  wire  _T_5192; // @[LoadQueue.scala 151:92:@5169.4]
  wire  _T_5193; // @[LoadQueue.scala 152:41:@5170.4]
  wire  _T_5194; // @[LoadQueue.scala 153:30:@5171.4]
  wire  conflict_1_4; // @[LoadQueue.scala 152:68:@5172.4]
  wire  _T_5196; // @[LoadQueue.scala 151:92:@5174.4]
  wire  _T_5197; // @[LoadQueue.scala 152:41:@5175.4]
  wire  _T_5198; // @[LoadQueue.scala 153:30:@5176.4]
  wire  conflict_1_5; // @[LoadQueue.scala 152:68:@5177.4]
  wire  _T_5200; // @[LoadQueue.scala 151:92:@5179.4]
  wire  _T_5201; // @[LoadQueue.scala 152:41:@5180.4]
  wire  _T_5202; // @[LoadQueue.scala 153:30:@5181.4]
  wire  conflict_1_6; // @[LoadQueue.scala 152:68:@5182.4]
  wire  _T_5204; // @[LoadQueue.scala 151:92:@5184.4]
  wire  _T_5205; // @[LoadQueue.scala 152:41:@5185.4]
  wire  _T_5206; // @[LoadQueue.scala 153:30:@5186.4]
  wire  conflict_1_7; // @[LoadQueue.scala 152:68:@5187.4]
  wire  _T_5208; // @[LoadQueue.scala 151:92:@5189.4]
  wire  _T_5209; // @[LoadQueue.scala 152:41:@5190.4]
  wire  _T_5210; // @[LoadQueue.scala 153:30:@5191.4]
  wire  conflict_2_0; // @[LoadQueue.scala 152:68:@5192.4]
  wire  _T_5212; // @[LoadQueue.scala 151:92:@5194.4]
  wire  _T_5213; // @[LoadQueue.scala 152:41:@5195.4]
  wire  _T_5214; // @[LoadQueue.scala 153:30:@5196.4]
  wire  conflict_2_1; // @[LoadQueue.scala 152:68:@5197.4]
  wire  _T_5216; // @[LoadQueue.scala 151:92:@5199.4]
  wire  _T_5217; // @[LoadQueue.scala 152:41:@5200.4]
  wire  _T_5218; // @[LoadQueue.scala 153:30:@5201.4]
  wire  conflict_2_2; // @[LoadQueue.scala 152:68:@5202.4]
  wire  _T_5220; // @[LoadQueue.scala 151:92:@5204.4]
  wire  _T_5221; // @[LoadQueue.scala 152:41:@5205.4]
  wire  _T_5222; // @[LoadQueue.scala 153:30:@5206.4]
  wire  conflict_2_3; // @[LoadQueue.scala 152:68:@5207.4]
  wire  _T_5224; // @[LoadQueue.scala 151:92:@5209.4]
  wire  _T_5225; // @[LoadQueue.scala 152:41:@5210.4]
  wire  _T_5226; // @[LoadQueue.scala 153:30:@5211.4]
  wire  conflict_2_4; // @[LoadQueue.scala 152:68:@5212.4]
  wire  _T_5228; // @[LoadQueue.scala 151:92:@5214.4]
  wire  _T_5229; // @[LoadQueue.scala 152:41:@5215.4]
  wire  _T_5230; // @[LoadQueue.scala 153:30:@5216.4]
  wire  conflict_2_5; // @[LoadQueue.scala 152:68:@5217.4]
  wire  _T_5232; // @[LoadQueue.scala 151:92:@5219.4]
  wire  _T_5233; // @[LoadQueue.scala 152:41:@5220.4]
  wire  _T_5234; // @[LoadQueue.scala 153:30:@5221.4]
  wire  conflict_2_6; // @[LoadQueue.scala 152:68:@5222.4]
  wire  _T_5236; // @[LoadQueue.scala 151:92:@5224.4]
  wire  _T_5237; // @[LoadQueue.scala 152:41:@5225.4]
  wire  _T_5238; // @[LoadQueue.scala 153:30:@5226.4]
  wire  conflict_2_7; // @[LoadQueue.scala 152:68:@5227.4]
  wire  _T_5240; // @[LoadQueue.scala 151:92:@5229.4]
  wire  _T_5241; // @[LoadQueue.scala 152:41:@5230.4]
  wire  _T_5242; // @[LoadQueue.scala 153:30:@5231.4]
  wire  conflict_3_0; // @[LoadQueue.scala 152:68:@5232.4]
  wire  _T_5244; // @[LoadQueue.scala 151:92:@5234.4]
  wire  _T_5245; // @[LoadQueue.scala 152:41:@5235.4]
  wire  _T_5246; // @[LoadQueue.scala 153:30:@5236.4]
  wire  conflict_3_1; // @[LoadQueue.scala 152:68:@5237.4]
  wire  _T_5248; // @[LoadQueue.scala 151:92:@5239.4]
  wire  _T_5249; // @[LoadQueue.scala 152:41:@5240.4]
  wire  _T_5250; // @[LoadQueue.scala 153:30:@5241.4]
  wire  conflict_3_2; // @[LoadQueue.scala 152:68:@5242.4]
  wire  _T_5252; // @[LoadQueue.scala 151:92:@5244.4]
  wire  _T_5253; // @[LoadQueue.scala 152:41:@5245.4]
  wire  _T_5254; // @[LoadQueue.scala 153:30:@5246.4]
  wire  conflict_3_3; // @[LoadQueue.scala 152:68:@5247.4]
  wire  _T_5256; // @[LoadQueue.scala 151:92:@5249.4]
  wire  _T_5257; // @[LoadQueue.scala 152:41:@5250.4]
  wire  _T_5258; // @[LoadQueue.scala 153:30:@5251.4]
  wire  conflict_3_4; // @[LoadQueue.scala 152:68:@5252.4]
  wire  _T_5260; // @[LoadQueue.scala 151:92:@5254.4]
  wire  _T_5261; // @[LoadQueue.scala 152:41:@5255.4]
  wire  _T_5262; // @[LoadQueue.scala 153:30:@5256.4]
  wire  conflict_3_5; // @[LoadQueue.scala 152:68:@5257.4]
  wire  _T_5264; // @[LoadQueue.scala 151:92:@5259.4]
  wire  _T_5265; // @[LoadQueue.scala 152:41:@5260.4]
  wire  _T_5266; // @[LoadQueue.scala 153:30:@5261.4]
  wire  conflict_3_6; // @[LoadQueue.scala 152:68:@5262.4]
  wire  _T_5268; // @[LoadQueue.scala 151:92:@5264.4]
  wire  _T_5269; // @[LoadQueue.scala 152:41:@5265.4]
  wire  _T_5270; // @[LoadQueue.scala 153:30:@5266.4]
  wire  conflict_3_7; // @[LoadQueue.scala 152:68:@5267.4]
  wire  _T_5272; // @[LoadQueue.scala 151:92:@5269.4]
  wire  _T_5273; // @[LoadQueue.scala 152:41:@5270.4]
  wire  _T_5274; // @[LoadQueue.scala 153:30:@5271.4]
  wire  conflict_4_0; // @[LoadQueue.scala 152:68:@5272.4]
  wire  _T_5276; // @[LoadQueue.scala 151:92:@5274.4]
  wire  _T_5277; // @[LoadQueue.scala 152:41:@5275.4]
  wire  _T_5278; // @[LoadQueue.scala 153:30:@5276.4]
  wire  conflict_4_1; // @[LoadQueue.scala 152:68:@5277.4]
  wire  _T_5280; // @[LoadQueue.scala 151:92:@5279.4]
  wire  _T_5281; // @[LoadQueue.scala 152:41:@5280.4]
  wire  _T_5282; // @[LoadQueue.scala 153:30:@5281.4]
  wire  conflict_4_2; // @[LoadQueue.scala 152:68:@5282.4]
  wire  _T_5284; // @[LoadQueue.scala 151:92:@5284.4]
  wire  _T_5285; // @[LoadQueue.scala 152:41:@5285.4]
  wire  _T_5286; // @[LoadQueue.scala 153:30:@5286.4]
  wire  conflict_4_3; // @[LoadQueue.scala 152:68:@5287.4]
  wire  _T_5288; // @[LoadQueue.scala 151:92:@5289.4]
  wire  _T_5289; // @[LoadQueue.scala 152:41:@5290.4]
  wire  _T_5290; // @[LoadQueue.scala 153:30:@5291.4]
  wire  conflict_4_4; // @[LoadQueue.scala 152:68:@5292.4]
  wire  _T_5292; // @[LoadQueue.scala 151:92:@5294.4]
  wire  _T_5293; // @[LoadQueue.scala 152:41:@5295.4]
  wire  _T_5294; // @[LoadQueue.scala 153:30:@5296.4]
  wire  conflict_4_5; // @[LoadQueue.scala 152:68:@5297.4]
  wire  _T_5296; // @[LoadQueue.scala 151:92:@5299.4]
  wire  _T_5297; // @[LoadQueue.scala 152:41:@5300.4]
  wire  _T_5298; // @[LoadQueue.scala 153:30:@5301.4]
  wire  conflict_4_6; // @[LoadQueue.scala 152:68:@5302.4]
  wire  _T_5300; // @[LoadQueue.scala 151:92:@5304.4]
  wire  _T_5301; // @[LoadQueue.scala 152:41:@5305.4]
  wire  _T_5302; // @[LoadQueue.scala 153:30:@5306.4]
  wire  conflict_4_7; // @[LoadQueue.scala 152:68:@5307.4]
  wire  _T_5304; // @[LoadQueue.scala 151:92:@5309.4]
  wire  _T_5305; // @[LoadQueue.scala 152:41:@5310.4]
  wire  _T_5306; // @[LoadQueue.scala 153:30:@5311.4]
  wire  conflict_5_0; // @[LoadQueue.scala 152:68:@5312.4]
  wire  _T_5308; // @[LoadQueue.scala 151:92:@5314.4]
  wire  _T_5309; // @[LoadQueue.scala 152:41:@5315.4]
  wire  _T_5310; // @[LoadQueue.scala 153:30:@5316.4]
  wire  conflict_5_1; // @[LoadQueue.scala 152:68:@5317.4]
  wire  _T_5312; // @[LoadQueue.scala 151:92:@5319.4]
  wire  _T_5313; // @[LoadQueue.scala 152:41:@5320.4]
  wire  _T_5314; // @[LoadQueue.scala 153:30:@5321.4]
  wire  conflict_5_2; // @[LoadQueue.scala 152:68:@5322.4]
  wire  _T_5316; // @[LoadQueue.scala 151:92:@5324.4]
  wire  _T_5317; // @[LoadQueue.scala 152:41:@5325.4]
  wire  _T_5318; // @[LoadQueue.scala 153:30:@5326.4]
  wire  conflict_5_3; // @[LoadQueue.scala 152:68:@5327.4]
  wire  _T_5320; // @[LoadQueue.scala 151:92:@5329.4]
  wire  _T_5321; // @[LoadQueue.scala 152:41:@5330.4]
  wire  _T_5322; // @[LoadQueue.scala 153:30:@5331.4]
  wire  conflict_5_4; // @[LoadQueue.scala 152:68:@5332.4]
  wire  _T_5324; // @[LoadQueue.scala 151:92:@5334.4]
  wire  _T_5325; // @[LoadQueue.scala 152:41:@5335.4]
  wire  _T_5326; // @[LoadQueue.scala 153:30:@5336.4]
  wire  conflict_5_5; // @[LoadQueue.scala 152:68:@5337.4]
  wire  _T_5328; // @[LoadQueue.scala 151:92:@5339.4]
  wire  _T_5329; // @[LoadQueue.scala 152:41:@5340.4]
  wire  _T_5330; // @[LoadQueue.scala 153:30:@5341.4]
  wire  conflict_5_6; // @[LoadQueue.scala 152:68:@5342.4]
  wire  _T_5332; // @[LoadQueue.scala 151:92:@5344.4]
  wire  _T_5333; // @[LoadQueue.scala 152:41:@5345.4]
  wire  _T_5334; // @[LoadQueue.scala 153:30:@5346.4]
  wire  conflict_5_7; // @[LoadQueue.scala 152:68:@5347.4]
  wire  _T_5336; // @[LoadQueue.scala 151:92:@5349.4]
  wire  _T_5337; // @[LoadQueue.scala 152:41:@5350.4]
  wire  _T_5338; // @[LoadQueue.scala 153:30:@5351.4]
  wire  conflict_6_0; // @[LoadQueue.scala 152:68:@5352.4]
  wire  _T_5340; // @[LoadQueue.scala 151:92:@5354.4]
  wire  _T_5341; // @[LoadQueue.scala 152:41:@5355.4]
  wire  _T_5342; // @[LoadQueue.scala 153:30:@5356.4]
  wire  conflict_6_1; // @[LoadQueue.scala 152:68:@5357.4]
  wire  _T_5344; // @[LoadQueue.scala 151:92:@5359.4]
  wire  _T_5345; // @[LoadQueue.scala 152:41:@5360.4]
  wire  _T_5346; // @[LoadQueue.scala 153:30:@5361.4]
  wire  conflict_6_2; // @[LoadQueue.scala 152:68:@5362.4]
  wire  _T_5348; // @[LoadQueue.scala 151:92:@5364.4]
  wire  _T_5349; // @[LoadQueue.scala 152:41:@5365.4]
  wire  _T_5350; // @[LoadQueue.scala 153:30:@5366.4]
  wire  conflict_6_3; // @[LoadQueue.scala 152:68:@5367.4]
  wire  _T_5352; // @[LoadQueue.scala 151:92:@5369.4]
  wire  _T_5353; // @[LoadQueue.scala 152:41:@5370.4]
  wire  _T_5354; // @[LoadQueue.scala 153:30:@5371.4]
  wire  conflict_6_4; // @[LoadQueue.scala 152:68:@5372.4]
  wire  _T_5356; // @[LoadQueue.scala 151:92:@5374.4]
  wire  _T_5357; // @[LoadQueue.scala 152:41:@5375.4]
  wire  _T_5358; // @[LoadQueue.scala 153:30:@5376.4]
  wire  conflict_6_5; // @[LoadQueue.scala 152:68:@5377.4]
  wire  _T_5360; // @[LoadQueue.scala 151:92:@5379.4]
  wire  _T_5361; // @[LoadQueue.scala 152:41:@5380.4]
  wire  _T_5362; // @[LoadQueue.scala 153:30:@5381.4]
  wire  conflict_6_6; // @[LoadQueue.scala 152:68:@5382.4]
  wire  _T_5364; // @[LoadQueue.scala 151:92:@5384.4]
  wire  _T_5365; // @[LoadQueue.scala 152:41:@5385.4]
  wire  _T_5366; // @[LoadQueue.scala 153:30:@5386.4]
  wire  conflict_6_7; // @[LoadQueue.scala 152:68:@5387.4]
  wire  _T_5368; // @[LoadQueue.scala 151:92:@5389.4]
  wire  _T_5369; // @[LoadQueue.scala 152:41:@5390.4]
  wire  _T_5370; // @[LoadQueue.scala 153:30:@5391.4]
  wire  conflict_7_0; // @[LoadQueue.scala 152:68:@5392.4]
  wire  _T_5372; // @[LoadQueue.scala 151:92:@5394.4]
  wire  _T_5373; // @[LoadQueue.scala 152:41:@5395.4]
  wire  _T_5374; // @[LoadQueue.scala 153:30:@5396.4]
  wire  conflict_7_1; // @[LoadQueue.scala 152:68:@5397.4]
  wire  _T_5376; // @[LoadQueue.scala 151:92:@5399.4]
  wire  _T_5377; // @[LoadQueue.scala 152:41:@5400.4]
  wire  _T_5378; // @[LoadQueue.scala 153:30:@5401.4]
  wire  conflict_7_2; // @[LoadQueue.scala 152:68:@5402.4]
  wire  _T_5380; // @[LoadQueue.scala 151:92:@5404.4]
  wire  _T_5381; // @[LoadQueue.scala 152:41:@5405.4]
  wire  _T_5382; // @[LoadQueue.scala 153:30:@5406.4]
  wire  conflict_7_3; // @[LoadQueue.scala 152:68:@5407.4]
  wire  _T_5384; // @[LoadQueue.scala 151:92:@5409.4]
  wire  _T_5385; // @[LoadQueue.scala 152:41:@5410.4]
  wire  _T_5386; // @[LoadQueue.scala 153:30:@5411.4]
  wire  conflict_7_4; // @[LoadQueue.scala 152:68:@5412.4]
  wire  _T_5388; // @[LoadQueue.scala 151:92:@5414.4]
  wire  _T_5389; // @[LoadQueue.scala 152:41:@5415.4]
  wire  _T_5390; // @[LoadQueue.scala 153:30:@5416.4]
  wire  conflict_7_5; // @[LoadQueue.scala 152:68:@5417.4]
  wire  _T_5392; // @[LoadQueue.scala 151:92:@5419.4]
  wire  _T_5393; // @[LoadQueue.scala 152:41:@5420.4]
  wire  _T_5394; // @[LoadQueue.scala 153:30:@5421.4]
  wire  conflict_7_6; // @[LoadQueue.scala 152:68:@5422.4]
  wire  _T_5396; // @[LoadQueue.scala 151:92:@5424.4]
  wire  _T_5397; // @[LoadQueue.scala 152:41:@5425.4]
  wire  _T_5398; // @[LoadQueue.scala 153:30:@5426.4]
  wire  conflict_7_7; // @[LoadQueue.scala 152:68:@5427.4]
  wire  _T_5767; // @[LoadQueue.scala 163:13:@5430.4]
  wire  storeAddrNotKnownFlags_0_0; // @[LoadQueue.scala 163:19:@5431.4]
  wire  _T_5770; // @[LoadQueue.scala 163:13:@5432.4]
  wire  storeAddrNotKnownFlags_0_1; // @[LoadQueue.scala 163:19:@5433.4]
  wire  _T_5773; // @[LoadQueue.scala 163:13:@5434.4]
  wire  storeAddrNotKnownFlags_0_2; // @[LoadQueue.scala 163:19:@5435.4]
  wire  _T_5776; // @[LoadQueue.scala 163:13:@5436.4]
  wire  storeAddrNotKnownFlags_0_3; // @[LoadQueue.scala 163:19:@5437.4]
  wire  _T_5779; // @[LoadQueue.scala 163:13:@5438.4]
  wire  storeAddrNotKnownFlags_0_4; // @[LoadQueue.scala 163:19:@5439.4]
  wire  _T_5782; // @[LoadQueue.scala 163:13:@5440.4]
  wire  storeAddrNotKnownFlags_0_5; // @[LoadQueue.scala 163:19:@5441.4]
  wire  _T_5785; // @[LoadQueue.scala 163:13:@5442.4]
  wire  storeAddrNotKnownFlags_0_6; // @[LoadQueue.scala 163:19:@5443.4]
  wire  _T_5788; // @[LoadQueue.scala 163:13:@5444.4]
  wire  storeAddrNotKnownFlags_0_7; // @[LoadQueue.scala 163:19:@5445.4]
  wire  storeAddrNotKnownFlags_1_0; // @[LoadQueue.scala 163:19:@5455.4]
  wire  storeAddrNotKnownFlags_1_1; // @[LoadQueue.scala 163:19:@5457.4]
  wire  storeAddrNotKnownFlags_1_2; // @[LoadQueue.scala 163:19:@5459.4]
  wire  storeAddrNotKnownFlags_1_3; // @[LoadQueue.scala 163:19:@5461.4]
  wire  storeAddrNotKnownFlags_1_4; // @[LoadQueue.scala 163:19:@5463.4]
  wire  storeAddrNotKnownFlags_1_5; // @[LoadQueue.scala 163:19:@5465.4]
  wire  storeAddrNotKnownFlags_1_6; // @[LoadQueue.scala 163:19:@5467.4]
  wire  storeAddrNotKnownFlags_1_7; // @[LoadQueue.scala 163:19:@5469.4]
  wire  storeAddrNotKnownFlags_2_0; // @[LoadQueue.scala 163:19:@5479.4]
  wire  storeAddrNotKnownFlags_2_1; // @[LoadQueue.scala 163:19:@5481.4]
  wire  storeAddrNotKnownFlags_2_2; // @[LoadQueue.scala 163:19:@5483.4]
  wire  storeAddrNotKnownFlags_2_3; // @[LoadQueue.scala 163:19:@5485.4]
  wire  storeAddrNotKnownFlags_2_4; // @[LoadQueue.scala 163:19:@5487.4]
  wire  storeAddrNotKnownFlags_2_5; // @[LoadQueue.scala 163:19:@5489.4]
  wire  storeAddrNotKnownFlags_2_6; // @[LoadQueue.scala 163:19:@5491.4]
  wire  storeAddrNotKnownFlags_2_7; // @[LoadQueue.scala 163:19:@5493.4]
  wire  storeAddrNotKnownFlags_3_0; // @[LoadQueue.scala 163:19:@5503.4]
  wire  storeAddrNotKnownFlags_3_1; // @[LoadQueue.scala 163:19:@5505.4]
  wire  storeAddrNotKnownFlags_3_2; // @[LoadQueue.scala 163:19:@5507.4]
  wire  storeAddrNotKnownFlags_3_3; // @[LoadQueue.scala 163:19:@5509.4]
  wire  storeAddrNotKnownFlags_3_4; // @[LoadQueue.scala 163:19:@5511.4]
  wire  storeAddrNotKnownFlags_3_5; // @[LoadQueue.scala 163:19:@5513.4]
  wire  storeAddrNotKnownFlags_3_6; // @[LoadQueue.scala 163:19:@5515.4]
  wire  storeAddrNotKnownFlags_3_7; // @[LoadQueue.scala 163:19:@5517.4]
  wire  storeAddrNotKnownFlags_4_0; // @[LoadQueue.scala 163:19:@5527.4]
  wire  storeAddrNotKnownFlags_4_1; // @[LoadQueue.scala 163:19:@5529.4]
  wire  storeAddrNotKnownFlags_4_2; // @[LoadQueue.scala 163:19:@5531.4]
  wire  storeAddrNotKnownFlags_4_3; // @[LoadQueue.scala 163:19:@5533.4]
  wire  storeAddrNotKnownFlags_4_4; // @[LoadQueue.scala 163:19:@5535.4]
  wire  storeAddrNotKnownFlags_4_5; // @[LoadQueue.scala 163:19:@5537.4]
  wire  storeAddrNotKnownFlags_4_6; // @[LoadQueue.scala 163:19:@5539.4]
  wire  storeAddrNotKnownFlags_4_7; // @[LoadQueue.scala 163:19:@5541.4]
  wire  storeAddrNotKnownFlags_5_0; // @[LoadQueue.scala 163:19:@5551.4]
  wire  storeAddrNotKnownFlags_5_1; // @[LoadQueue.scala 163:19:@5553.4]
  wire  storeAddrNotKnownFlags_5_2; // @[LoadQueue.scala 163:19:@5555.4]
  wire  storeAddrNotKnownFlags_5_3; // @[LoadQueue.scala 163:19:@5557.4]
  wire  storeAddrNotKnownFlags_5_4; // @[LoadQueue.scala 163:19:@5559.4]
  wire  storeAddrNotKnownFlags_5_5; // @[LoadQueue.scala 163:19:@5561.4]
  wire  storeAddrNotKnownFlags_5_6; // @[LoadQueue.scala 163:19:@5563.4]
  wire  storeAddrNotKnownFlags_5_7; // @[LoadQueue.scala 163:19:@5565.4]
  wire  storeAddrNotKnownFlags_6_0; // @[LoadQueue.scala 163:19:@5575.4]
  wire  storeAddrNotKnownFlags_6_1; // @[LoadQueue.scala 163:19:@5577.4]
  wire  storeAddrNotKnownFlags_6_2; // @[LoadQueue.scala 163:19:@5579.4]
  wire  storeAddrNotKnownFlags_6_3; // @[LoadQueue.scala 163:19:@5581.4]
  wire  storeAddrNotKnownFlags_6_4; // @[LoadQueue.scala 163:19:@5583.4]
  wire  storeAddrNotKnownFlags_6_5; // @[LoadQueue.scala 163:19:@5585.4]
  wire  storeAddrNotKnownFlags_6_6; // @[LoadQueue.scala 163:19:@5587.4]
  wire  storeAddrNotKnownFlags_6_7; // @[LoadQueue.scala 163:19:@5589.4]
  wire  storeAddrNotKnownFlags_7_0; // @[LoadQueue.scala 163:19:@5599.4]
  wire  storeAddrNotKnownFlags_7_1; // @[LoadQueue.scala 163:19:@5601.4]
  wire  storeAddrNotKnownFlags_7_2; // @[LoadQueue.scala 163:19:@5603.4]
  wire  storeAddrNotKnownFlags_7_3; // @[LoadQueue.scala 163:19:@5605.4]
  wire  storeAddrNotKnownFlags_7_4; // @[LoadQueue.scala 163:19:@5607.4]
  wire  storeAddrNotKnownFlags_7_5; // @[LoadQueue.scala 163:19:@5609.4]
  wire  storeAddrNotKnownFlags_7_6; // @[LoadQueue.scala 163:19:@5611.4]
  wire  storeAddrNotKnownFlags_7_7; // @[LoadQueue.scala 163:19:@5613.4]
  wire [7:0] _T_6122; // @[Mux.scala 19:72:@5720.4]
  wire [7:0] _T_6124; // @[Mux.scala 19:72:@5721.4]
  wire [7:0] _T_6131; // @[Mux.scala 19:72:@5728.4]
  wire [7:0] _T_6133; // @[Mux.scala 19:72:@5729.4]
  wire [7:0] _T_6140; // @[Mux.scala 19:72:@5736.4]
  wire [7:0] _T_6142; // @[Mux.scala 19:72:@5737.4]
  wire [7:0] _T_6149; // @[Mux.scala 19:72:@5744.4]
  wire [7:0] _T_6151; // @[Mux.scala 19:72:@5745.4]
  wire [7:0] _T_6158; // @[Mux.scala 19:72:@5752.4]
  wire [7:0] _T_6160; // @[Mux.scala 19:72:@5753.4]
  wire [7:0] _T_6167; // @[Mux.scala 19:72:@5760.4]
  wire [7:0] _T_6169; // @[Mux.scala 19:72:@5761.4]
  wire [7:0] _T_6176; // @[Mux.scala 19:72:@5768.4]
  wire [7:0] _T_6178; // @[Mux.scala 19:72:@5769.4]
  wire [7:0] _T_6185; // @[Mux.scala 19:72:@5776.4]
  wire [7:0] _T_6187; // @[Mux.scala 19:72:@5777.4]
  wire [7:0] _T_6188; // @[Mux.scala 19:72:@5778.4]
  wire [7:0] _T_6189; // @[Mux.scala 19:72:@5779.4]
  wire [7:0] _T_6190; // @[Mux.scala 19:72:@5780.4]
  wire [7:0] _T_6191; // @[Mux.scala 19:72:@5781.4]
  wire [7:0] _T_6192; // @[Mux.scala 19:72:@5782.4]
  wire [7:0] _T_6193; // @[Mux.scala 19:72:@5783.4]
  wire [7:0] _T_6194; // @[Mux.scala 19:72:@5784.4]
  wire [7:0] _T_6436; // @[Mux.scala 19:72:@5902.4]
  wire [7:0] _T_6438; // @[Mux.scala 19:72:@5903.4]
  wire [7:0] _T_6445; // @[Mux.scala 19:72:@5910.4]
  wire [7:0] _T_6447; // @[Mux.scala 19:72:@5911.4]
  wire [7:0] _T_6454; // @[Mux.scala 19:72:@5918.4]
  wire [7:0] _T_6456; // @[Mux.scala 19:72:@5919.4]
  wire [7:0] _T_6463; // @[Mux.scala 19:72:@5926.4]
  wire [7:0] _T_6465; // @[Mux.scala 19:72:@5927.4]
  wire [7:0] _T_6472; // @[Mux.scala 19:72:@5934.4]
  wire [7:0] _T_6474; // @[Mux.scala 19:72:@5935.4]
  wire [7:0] _T_6481; // @[Mux.scala 19:72:@5942.4]
  wire [7:0] _T_6483; // @[Mux.scala 19:72:@5943.4]
  wire [7:0] _T_6490; // @[Mux.scala 19:72:@5950.4]
  wire [7:0] _T_6492; // @[Mux.scala 19:72:@5951.4]
  wire [7:0] _T_6499; // @[Mux.scala 19:72:@5958.4]
  wire [7:0] _T_6501; // @[Mux.scala 19:72:@5959.4]
  wire [7:0] _T_6502; // @[Mux.scala 19:72:@5960.4]
  wire [7:0] _T_6503; // @[Mux.scala 19:72:@5961.4]
  wire [7:0] _T_6504; // @[Mux.scala 19:72:@5962.4]
  wire [7:0] _T_6505; // @[Mux.scala 19:72:@5963.4]
  wire [7:0] _T_6506; // @[Mux.scala 19:72:@5964.4]
  wire [7:0] _T_6507; // @[Mux.scala 19:72:@5965.4]
  wire [7:0] _T_6508; // @[Mux.scala 19:72:@5966.4]
  wire [7:0] _T_6750; // @[Mux.scala 19:72:@6084.4]
  wire [7:0] _T_6752; // @[Mux.scala 19:72:@6085.4]
  wire [7:0] _T_6759; // @[Mux.scala 19:72:@6092.4]
  wire [7:0] _T_6761; // @[Mux.scala 19:72:@6093.4]
  wire [7:0] _T_6768; // @[Mux.scala 19:72:@6100.4]
  wire [7:0] _T_6770; // @[Mux.scala 19:72:@6101.4]
  wire [7:0] _T_6777; // @[Mux.scala 19:72:@6108.4]
  wire [7:0] _T_6779; // @[Mux.scala 19:72:@6109.4]
  wire [7:0] _T_6786; // @[Mux.scala 19:72:@6116.4]
  wire [7:0] _T_6788; // @[Mux.scala 19:72:@6117.4]
  wire [7:0] _T_6795; // @[Mux.scala 19:72:@6124.4]
  wire [7:0] _T_6797; // @[Mux.scala 19:72:@6125.4]
  wire [7:0] _T_6804; // @[Mux.scala 19:72:@6132.4]
  wire [7:0] _T_6806; // @[Mux.scala 19:72:@6133.4]
  wire [7:0] _T_6813; // @[Mux.scala 19:72:@6140.4]
  wire [7:0] _T_6815; // @[Mux.scala 19:72:@6141.4]
  wire [7:0] _T_6816; // @[Mux.scala 19:72:@6142.4]
  wire [7:0] _T_6817; // @[Mux.scala 19:72:@6143.4]
  wire [7:0] _T_6818; // @[Mux.scala 19:72:@6144.4]
  wire [7:0] _T_6819; // @[Mux.scala 19:72:@6145.4]
  wire [7:0] _T_6820; // @[Mux.scala 19:72:@6146.4]
  wire [7:0] _T_6821; // @[Mux.scala 19:72:@6147.4]
  wire [7:0] _T_6822; // @[Mux.scala 19:72:@6148.4]
  wire [7:0] _T_7064; // @[Mux.scala 19:72:@6266.4]
  wire [7:0] _T_7066; // @[Mux.scala 19:72:@6267.4]
  wire [7:0] _T_7073; // @[Mux.scala 19:72:@6274.4]
  wire [7:0] _T_7075; // @[Mux.scala 19:72:@6275.4]
  wire [7:0] _T_7082; // @[Mux.scala 19:72:@6282.4]
  wire [7:0] _T_7084; // @[Mux.scala 19:72:@6283.4]
  wire [7:0] _T_7091; // @[Mux.scala 19:72:@6290.4]
  wire [7:0] _T_7093; // @[Mux.scala 19:72:@6291.4]
  wire [7:0] _T_7100; // @[Mux.scala 19:72:@6298.4]
  wire [7:0] _T_7102; // @[Mux.scala 19:72:@6299.4]
  wire [7:0] _T_7109; // @[Mux.scala 19:72:@6306.4]
  wire [7:0] _T_7111; // @[Mux.scala 19:72:@6307.4]
  wire [7:0] _T_7118; // @[Mux.scala 19:72:@6314.4]
  wire [7:0] _T_7120; // @[Mux.scala 19:72:@6315.4]
  wire [7:0] _T_7127; // @[Mux.scala 19:72:@6322.4]
  wire [7:0] _T_7129; // @[Mux.scala 19:72:@6323.4]
  wire [7:0] _T_7130; // @[Mux.scala 19:72:@6324.4]
  wire [7:0] _T_7131; // @[Mux.scala 19:72:@6325.4]
  wire [7:0] _T_7132; // @[Mux.scala 19:72:@6326.4]
  wire [7:0] _T_7133; // @[Mux.scala 19:72:@6327.4]
  wire [7:0] _T_7134; // @[Mux.scala 19:72:@6328.4]
  wire [7:0] _T_7135; // @[Mux.scala 19:72:@6329.4]
  wire [7:0] _T_7136; // @[Mux.scala 19:72:@6330.4]
  wire [7:0] _T_7378; // @[Mux.scala 19:72:@6448.4]
  wire [7:0] _T_7380; // @[Mux.scala 19:72:@6449.4]
  wire [7:0] _T_7387; // @[Mux.scala 19:72:@6456.4]
  wire [7:0] _T_7389; // @[Mux.scala 19:72:@6457.4]
  wire [7:0] _T_7396; // @[Mux.scala 19:72:@6464.4]
  wire [7:0] _T_7398; // @[Mux.scala 19:72:@6465.4]
  wire [7:0] _T_7405; // @[Mux.scala 19:72:@6472.4]
  wire [7:0] _T_7407; // @[Mux.scala 19:72:@6473.4]
  wire [7:0] _T_7414; // @[Mux.scala 19:72:@6480.4]
  wire [7:0] _T_7416; // @[Mux.scala 19:72:@6481.4]
  wire [7:0] _T_7423; // @[Mux.scala 19:72:@6488.4]
  wire [7:0] _T_7425; // @[Mux.scala 19:72:@6489.4]
  wire [7:0] _T_7432; // @[Mux.scala 19:72:@6496.4]
  wire [7:0] _T_7434; // @[Mux.scala 19:72:@6497.4]
  wire [7:0] _T_7441; // @[Mux.scala 19:72:@6504.4]
  wire [7:0] _T_7443; // @[Mux.scala 19:72:@6505.4]
  wire [7:0] _T_7444; // @[Mux.scala 19:72:@6506.4]
  wire [7:0] _T_7445; // @[Mux.scala 19:72:@6507.4]
  wire [7:0] _T_7446; // @[Mux.scala 19:72:@6508.4]
  wire [7:0] _T_7447; // @[Mux.scala 19:72:@6509.4]
  wire [7:0] _T_7448; // @[Mux.scala 19:72:@6510.4]
  wire [7:0] _T_7449; // @[Mux.scala 19:72:@6511.4]
  wire [7:0] _T_7450; // @[Mux.scala 19:72:@6512.4]
  wire [7:0] _T_7692; // @[Mux.scala 19:72:@6630.4]
  wire [7:0] _T_7694; // @[Mux.scala 19:72:@6631.4]
  wire [7:0] _T_7701; // @[Mux.scala 19:72:@6638.4]
  wire [7:0] _T_7703; // @[Mux.scala 19:72:@6639.4]
  wire [7:0] _T_7710; // @[Mux.scala 19:72:@6646.4]
  wire [7:0] _T_7712; // @[Mux.scala 19:72:@6647.4]
  wire [7:0] _T_7719; // @[Mux.scala 19:72:@6654.4]
  wire [7:0] _T_7721; // @[Mux.scala 19:72:@6655.4]
  wire [7:0] _T_7728; // @[Mux.scala 19:72:@6662.4]
  wire [7:0] _T_7730; // @[Mux.scala 19:72:@6663.4]
  wire [7:0] _T_7737; // @[Mux.scala 19:72:@6670.4]
  wire [7:0] _T_7739; // @[Mux.scala 19:72:@6671.4]
  wire [7:0] _T_7746; // @[Mux.scala 19:72:@6678.4]
  wire [7:0] _T_7748; // @[Mux.scala 19:72:@6679.4]
  wire [7:0] _T_7755; // @[Mux.scala 19:72:@6686.4]
  wire [7:0] _T_7757; // @[Mux.scala 19:72:@6687.4]
  wire [7:0] _T_7758; // @[Mux.scala 19:72:@6688.4]
  wire [7:0] _T_7759; // @[Mux.scala 19:72:@6689.4]
  wire [7:0] _T_7760; // @[Mux.scala 19:72:@6690.4]
  wire [7:0] _T_7761; // @[Mux.scala 19:72:@6691.4]
  wire [7:0] _T_7762; // @[Mux.scala 19:72:@6692.4]
  wire [7:0] _T_7763; // @[Mux.scala 19:72:@6693.4]
  wire [7:0] _T_7764; // @[Mux.scala 19:72:@6694.4]
  wire [7:0] _T_8006; // @[Mux.scala 19:72:@6812.4]
  wire [7:0] _T_8008; // @[Mux.scala 19:72:@6813.4]
  wire [7:0] _T_8015; // @[Mux.scala 19:72:@6820.4]
  wire [7:0] _T_8017; // @[Mux.scala 19:72:@6821.4]
  wire [7:0] _T_8024; // @[Mux.scala 19:72:@6828.4]
  wire [7:0] _T_8026; // @[Mux.scala 19:72:@6829.4]
  wire [7:0] _T_8033; // @[Mux.scala 19:72:@6836.4]
  wire [7:0] _T_8035; // @[Mux.scala 19:72:@6837.4]
  wire [7:0] _T_8042; // @[Mux.scala 19:72:@6844.4]
  wire [7:0] _T_8044; // @[Mux.scala 19:72:@6845.4]
  wire [7:0] _T_8051; // @[Mux.scala 19:72:@6852.4]
  wire [7:0] _T_8053; // @[Mux.scala 19:72:@6853.4]
  wire [7:0] _T_8060; // @[Mux.scala 19:72:@6860.4]
  wire [7:0] _T_8062; // @[Mux.scala 19:72:@6861.4]
  wire [7:0] _T_8069; // @[Mux.scala 19:72:@6868.4]
  wire [7:0] _T_8071; // @[Mux.scala 19:72:@6869.4]
  wire [7:0] _T_8072; // @[Mux.scala 19:72:@6870.4]
  wire [7:0] _T_8073; // @[Mux.scala 19:72:@6871.4]
  wire [7:0] _T_8074; // @[Mux.scala 19:72:@6872.4]
  wire [7:0] _T_8075; // @[Mux.scala 19:72:@6873.4]
  wire [7:0] _T_8076; // @[Mux.scala 19:72:@6874.4]
  wire [7:0] _T_8077; // @[Mux.scala 19:72:@6875.4]
  wire [7:0] _T_8078; // @[Mux.scala 19:72:@6876.4]
  wire [7:0] _T_8320; // @[Mux.scala 19:72:@6994.4]
  wire [7:0] _T_8322; // @[Mux.scala 19:72:@6995.4]
  wire [7:0] _T_8329; // @[Mux.scala 19:72:@7002.4]
  wire [7:0] _T_8331; // @[Mux.scala 19:72:@7003.4]
  wire [7:0] _T_8338; // @[Mux.scala 19:72:@7010.4]
  wire [7:0] _T_8340; // @[Mux.scala 19:72:@7011.4]
  wire [7:0] _T_8347; // @[Mux.scala 19:72:@7018.4]
  wire [7:0] _T_8349; // @[Mux.scala 19:72:@7019.4]
  wire [7:0] _T_8356; // @[Mux.scala 19:72:@7026.4]
  wire [7:0] _T_8358; // @[Mux.scala 19:72:@7027.4]
  wire [7:0] _T_8365; // @[Mux.scala 19:72:@7034.4]
  wire [7:0] _T_8367; // @[Mux.scala 19:72:@7035.4]
  wire [7:0] _T_8374; // @[Mux.scala 19:72:@7042.4]
  wire [7:0] _T_8376; // @[Mux.scala 19:72:@7043.4]
  wire [7:0] _T_8383; // @[Mux.scala 19:72:@7050.4]
  wire [7:0] _T_8385; // @[Mux.scala 19:72:@7051.4]
  wire [7:0] _T_8386; // @[Mux.scala 19:72:@7052.4]
  wire [7:0] _T_8387; // @[Mux.scala 19:72:@7053.4]
  wire [7:0] _T_8388; // @[Mux.scala 19:72:@7054.4]
  wire [7:0] _T_8389; // @[Mux.scala 19:72:@7055.4]
  wire [7:0] _T_8390; // @[Mux.scala 19:72:@7056.4]
  wire [7:0] _T_8391; // @[Mux.scala 19:72:@7057.4]
  wire [7:0] _T_8392; // @[Mux.scala 19:72:@7058.4]
  reg  conflictPReg_0_0; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_83;
  reg  conflictPReg_0_1; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_84;
  reg  conflictPReg_0_2; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_85;
  reg  conflictPReg_0_3; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_86;
  reg  conflictPReg_0_4; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_87;
  reg  conflictPReg_0_5; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_88;
  reg  conflictPReg_0_6; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_89;
  reg  conflictPReg_0_7; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_90;
  reg  conflictPReg_1_0; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_91;
  reg  conflictPReg_1_1; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_92;
  reg  conflictPReg_1_2; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_93;
  reg  conflictPReg_1_3; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_94;
  reg  conflictPReg_1_4; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_95;
  reg  conflictPReg_1_5; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_96;
  reg  conflictPReg_1_6; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_97;
  reg  conflictPReg_1_7; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_98;
  reg  conflictPReg_2_0; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_99;
  reg  conflictPReg_2_1; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_100;
  reg  conflictPReg_2_2; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_101;
  reg  conflictPReg_2_3; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_102;
  reg  conflictPReg_2_4; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_103;
  reg  conflictPReg_2_5; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_104;
  reg  conflictPReg_2_6; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_105;
  reg  conflictPReg_2_7; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_106;
  reg  conflictPReg_3_0; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_107;
  reg  conflictPReg_3_1; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_108;
  reg  conflictPReg_3_2; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_109;
  reg  conflictPReg_3_3; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_110;
  reg  conflictPReg_3_4; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_111;
  reg  conflictPReg_3_5; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_112;
  reg  conflictPReg_3_6; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_113;
  reg  conflictPReg_3_7; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_114;
  reg  conflictPReg_4_0; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_115;
  reg  conflictPReg_4_1; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_116;
  reg  conflictPReg_4_2; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_117;
  reg  conflictPReg_4_3; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_118;
  reg  conflictPReg_4_4; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_119;
  reg  conflictPReg_4_5; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_120;
  reg  conflictPReg_4_6; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_121;
  reg  conflictPReg_4_7; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_122;
  reg  conflictPReg_5_0; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_123;
  reg  conflictPReg_5_1; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_124;
  reg  conflictPReg_5_2; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_125;
  reg  conflictPReg_5_3; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_126;
  reg  conflictPReg_5_4; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_127;
  reg  conflictPReg_5_5; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_128;
  reg  conflictPReg_5_6; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_129;
  reg  conflictPReg_5_7; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_130;
  reg  conflictPReg_6_0; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_131;
  reg  conflictPReg_6_1; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_132;
  reg  conflictPReg_6_2; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_133;
  reg  conflictPReg_6_3; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_134;
  reg  conflictPReg_6_4; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_135;
  reg  conflictPReg_6_5; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_136;
  reg  conflictPReg_6_6; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_137;
  reg  conflictPReg_6_7; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_138;
  reg  conflictPReg_7_0; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_139;
  reg  conflictPReg_7_1; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_140;
  reg  conflictPReg_7_2; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_141;
  reg  conflictPReg_7_3; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_142;
  reg  conflictPReg_7_4; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_143;
  reg  conflictPReg_7_5; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_144;
  reg  conflictPReg_7_6; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_145;
  reg  conflictPReg_7_7; // @[LoadQueue.scala 166:29:@7143.4]
  reg [31:0] _RAND_146;
  wire [7:0] _T_14502; // @[Mux.scala 19:72:@7306.4]
  wire [7:0] _T_14504; // @[Mux.scala 19:72:@7307.4]
  wire [7:0] _T_14511; // @[Mux.scala 19:72:@7314.4]
  wire [7:0] _T_14513; // @[Mux.scala 19:72:@7315.4]
  wire [7:0] _T_14520; // @[Mux.scala 19:72:@7322.4]
  wire [7:0] _T_14522; // @[Mux.scala 19:72:@7323.4]
  wire [7:0] _T_14529; // @[Mux.scala 19:72:@7330.4]
  wire [7:0] _T_14531; // @[Mux.scala 19:72:@7331.4]
  wire [7:0] _T_14538; // @[Mux.scala 19:72:@7338.4]
  wire [7:0] _T_14540; // @[Mux.scala 19:72:@7339.4]
  wire [7:0] _T_14547; // @[Mux.scala 19:72:@7346.4]
  wire [7:0] _T_14549; // @[Mux.scala 19:72:@7347.4]
  wire [7:0] _T_14556; // @[Mux.scala 19:72:@7354.4]
  wire [7:0] _T_14558; // @[Mux.scala 19:72:@7355.4]
  wire [7:0] _T_14565; // @[Mux.scala 19:72:@7362.4]
  wire [7:0] _T_14567; // @[Mux.scala 19:72:@7363.4]
  wire [7:0] _T_14568; // @[Mux.scala 19:72:@7364.4]
  wire [7:0] _T_14569; // @[Mux.scala 19:72:@7365.4]
  wire [7:0] _T_14570; // @[Mux.scala 19:72:@7366.4]
  wire [7:0] _T_14571; // @[Mux.scala 19:72:@7367.4]
  wire [7:0] _T_14572; // @[Mux.scala 19:72:@7368.4]
  wire [7:0] _T_14573; // @[Mux.scala 19:72:@7369.4]
  wire [7:0] _T_14574; // @[Mux.scala 19:72:@7370.4]
  wire [7:0] _T_14816; // @[Mux.scala 19:72:@7488.4]
  wire [7:0] _T_14818; // @[Mux.scala 19:72:@7489.4]
  wire [7:0] _T_14825; // @[Mux.scala 19:72:@7496.4]
  wire [7:0] _T_14827; // @[Mux.scala 19:72:@7497.4]
  wire [7:0] _T_14834; // @[Mux.scala 19:72:@7504.4]
  wire [7:0] _T_14836; // @[Mux.scala 19:72:@7505.4]
  wire [7:0] _T_14843; // @[Mux.scala 19:72:@7512.4]
  wire [7:0] _T_14845; // @[Mux.scala 19:72:@7513.4]
  wire [7:0] _T_14852; // @[Mux.scala 19:72:@7520.4]
  wire [7:0] _T_14854; // @[Mux.scala 19:72:@7521.4]
  wire [7:0] _T_14861; // @[Mux.scala 19:72:@7528.4]
  wire [7:0] _T_14863; // @[Mux.scala 19:72:@7529.4]
  wire [7:0] _T_14870; // @[Mux.scala 19:72:@7536.4]
  wire [7:0] _T_14872; // @[Mux.scala 19:72:@7537.4]
  wire [7:0] _T_14879; // @[Mux.scala 19:72:@7544.4]
  wire [7:0] _T_14881; // @[Mux.scala 19:72:@7545.4]
  wire [7:0] _T_14882; // @[Mux.scala 19:72:@7546.4]
  wire [7:0] _T_14883; // @[Mux.scala 19:72:@7547.4]
  wire [7:0] _T_14884; // @[Mux.scala 19:72:@7548.4]
  wire [7:0] _T_14885; // @[Mux.scala 19:72:@7549.4]
  wire [7:0] _T_14886; // @[Mux.scala 19:72:@7550.4]
  wire [7:0] _T_14887; // @[Mux.scala 19:72:@7551.4]
  wire [7:0] _T_14888; // @[Mux.scala 19:72:@7552.4]
  wire [7:0] _T_15130; // @[Mux.scala 19:72:@7670.4]
  wire [7:0] _T_15132; // @[Mux.scala 19:72:@7671.4]
  wire [7:0] _T_15139; // @[Mux.scala 19:72:@7678.4]
  wire [7:0] _T_15141; // @[Mux.scala 19:72:@7679.4]
  wire [7:0] _T_15148; // @[Mux.scala 19:72:@7686.4]
  wire [7:0] _T_15150; // @[Mux.scala 19:72:@7687.4]
  wire [7:0] _T_15157; // @[Mux.scala 19:72:@7694.4]
  wire [7:0] _T_15159; // @[Mux.scala 19:72:@7695.4]
  wire [7:0] _T_15166; // @[Mux.scala 19:72:@7702.4]
  wire [7:0] _T_15168; // @[Mux.scala 19:72:@7703.4]
  wire [7:0] _T_15175; // @[Mux.scala 19:72:@7710.4]
  wire [7:0] _T_15177; // @[Mux.scala 19:72:@7711.4]
  wire [7:0] _T_15184; // @[Mux.scala 19:72:@7718.4]
  wire [7:0] _T_15186; // @[Mux.scala 19:72:@7719.4]
  wire [7:0] _T_15193; // @[Mux.scala 19:72:@7726.4]
  wire [7:0] _T_15195; // @[Mux.scala 19:72:@7727.4]
  wire [7:0] _T_15196; // @[Mux.scala 19:72:@7728.4]
  wire [7:0] _T_15197; // @[Mux.scala 19:72:@7729.4]
  wire [7:0] _T_15198; // @[Mux.scala 19:72:@7730.4]
  wire [7:0] _T_15199; // @[Mux.scala 19:72:@7731.4]
  wire [7:0] _T_15200; // @[Mux.scala 19:72:@7732.4]
  wire [7:0] _T_15201; // @[Mux.scala 19:72:@7733.4]
  wire [7:0] _T_15202; // @[Mux.scala 19:72:@7734.4]
  wire [7:0] _T_15444; // @[Mux.scala 19:72:@7852.4]
  wire [7:0] _T_15446; // @[Mux.scala 19:72:@7853.4]
  wire [7:0] _T_15453; // @[Mux.scala 19:72:@7860.4]
  wire [7:0] _T_15455; // @[Mux.scala 19:72:@7861.4]
  wire [7:0] _T_15462; // @[Mux.scala 19:72:@7868.4]
  wire [7:0] _T_15464; // @[Mux.scala 19:72:@7869.4]
  wire [7:0] _T_15471; // @[Mux.scala 19:72:@7876.4]
  wire [7:0] _T_15473; // @[Mux.scala 19:72:@7877.4]
  wire [7:0] _T_15480; // @[Mux.scala 19:72:@7884.4]
  wire [7:0] _T_15482; // @[Mux.scala 19:72:@7885.4]
  wire [7:0] _T_15489; // @[Mux.scala 19:72:@7892.4]
  wire [7:0] _T_15491; // @[Mux.scala 19:72:@7893.4]
  wire [7:0] _T_15498; // @[Mux.scala 19:72:@7900.4]
  wire [7:0] _T_15500; // @[Mux.scala 19:72:@7901.4]
  wire [7:0] _T_15507; // @[Mux.scala 19:72:@7908.4]
  wire [7:0] _T_15509; // @[Mux.scala 19:72:@7909.4]
  wire [7:0] _T_15510; // @[Mux.scala 19:72:@7910.4]
  wire [7:0] _T_15511; // @[Mux.scala 19:72:@7911.4]
  wire [7:0] _T_15512; // @[Mux.scala 19:72:@7912.4]
  wire [7:0] _T_15513; // @[Mux.scala 19:72:@7913.4]
  wire [7:0] _T_15514; // @[Mux.scala 19:72:@7914.4]
  wire [7:0] _T_15515; // @[Mux.scala 19:72:@7915.4]
  wire [7:0] _T_15516; // @[Mux.scala 19:72:@7916.4]
  wire [7:0] _T_15758; // @[Mux.scala 19:72:@8034.4]
  wire [7:0] _T_15760; // @[Mux.scala 19:72:@8035.4]
  wire [7:0] _T_15767; // @[Mux.scala 19:72:@8042.4]
  wire [7:0] _T_15769; // @[Mux.scala 19:72:@8043.4]
  wire [7:0] _T_15776; // @[Mux.scala 19:72:@8050.4]
  wire [7:0] _T_15778; // @[Mux.scala 19:72:@8051.4]
  wire [7:0] _T_15785; // @[Mux.scala 19:72:@8058.4]
  wire [7:0] _T_15787; // @[Mux.scala 19:72:@8059.4]
  wire [7:0] _T_15794; // @[Mux.scala 19:72:@8066.4]
  wire [7:0] _T_15796; // @[Mux.scala 19:72:@8067.4]
  wire [7:0] _T_15803; // @[Mux.scala 19:72:@8074.4]
  wire [7:0] _T_15805; // @[Mux.scala 19:72:@8075.4]
  wire [7:0] _T_15812; // @[Mux.scala 19:72:@8082.4]
  wire [7:0] _T_15814; // @[Mux.scala 19:72:@8083.4]
  wire [7:0] _T_15821; // @[Mux.scala 19:72:@8090.4]
  wire [7:0] _T_15823; // @[Mux.scala 19:72:@8091.4]
  wire [7:0] _T_15824; // @[Mux.scala 19:72:@8092.4]
  wire [7:0] _T_15825; // @[Mux.scala 19:72:@8093.4]
  wire [7:0] _T_15826; // @[Mux.scala 19:72:@8094.4]
  wire [7:0] _T_15827; // @[Mux.scala 19:72:@8095.4]
  wire [7:0] _T_15828; // @[Mux.scala 19:72:@8096.4]
  wire [7:0] _T_15829; // @[Mux.scala 19:72:@8097.4]
  wire [7:0] _T_15830; // @[Mux.scala 19:72:@8098.4]
  wire [7:0] _T_16072; // @[Mux.scala 19:72:@8216.4]
  wire [7:0] _T_16074; // @[Mux.scala 19:72:@8217.4]
  wire [7:0] _T_16081; // @[Mux.scala 19:72:@8224.4]
  wire [7:0] _T_16083; // @[Mux.scala 19:72:@8225.4]
  wire [7:0] _T_16090; // @[Mux.scala 19:72:@8232.4]
  wire [7:0] _T_16092; // @[Mux.scala 19:72:@8233.4]
  wire [7:0] _T_16099; // @[Mux.scala 19:72:@8240.4]
  wire [7:0] _T_16101; // @[Mux.scala 19:72:@8241.4]
  wire [7:0] _T_16108; // @[Mux.scala 19:72:@8248.4]
  wire [7:0] _T_16110; // @[Mux.scala 19:72:@8249.4]
  wire [7:0] _T_16117; // @[Mux.scala 19:72:@8256.4]
  wire [7:0] _T_16119; // @[Mux.scala 19:72:@8257.4]
  wire [7:0] _T_16126; // @[Mux.scala 19:72:@8264.4]
  wire [7:0] _T_16128; // @[Mux.scala 19:72:@8265.4]
  wire [7:0] _T_16135; // @[Mux.scala 19:72:@8272.4]
  wire [7:0] _T_16137; // @[Mux.scala 19:72:@8273.4]
  wire [7:0] _T_16138; // @[Mux.scala 19:72:@8274.4]
  wire [7:0] _T_16139; // @[Mux.scala 19:72:@8275.4]
  wire [7:0] _T_16140; // @[Mux.scala 19:72:@8276.4]
  wire [7:0] _T_16141; // @[Mux.scala 19:72:@8277.4]
  wire [7:0] _T_16142; // @[Mux.scala 19:72:@8278.4]
  wire [7:0] _T_16143; // @[Mux.scala 19:72:@8279.4]
  wire [7:0] _T_16144; // @[Mux.scala 19:72:@8280.4]
  wire [7:0] _T_16386; // @[Mux.scala 19:72:@8398.4]
  wire [7:0] _T_16388; // @[Mux.scala 19:72:@8399.4]
  wire [7:0] _T_16395; // @[Mux.scala 19:72:@8406.4]
  wire [7:0] _T_16397; // @[Mux.scala 19:72:@8407.4]
  wire [7:0] _T_16404; // @[Mux.scala 19:72:@8414.4]
  wire [7:0] _T_16406; // @[Mux.scala 19:72:@8415.4]
  wire [7:0] _T_16413; // @[Mux.scala 19:72:@8422.4]
  wire [7:0] _T_16415; // @[Mux.scala 19:72:@8423.4]
  wire [7:0] _T_16422; // @[Mux.scala 19:72:@8430.4]
  wire [7:0] _T_16424; // @[Mux.scala 19:72:@8431.4]
  wire [7:0] _T_16431; // @[Mux.scala 19:72:@8438.4]
  wire [7:0] _T_16433; // @[Mux.scala 19:72:@8439.4]
  wire [7:0] _T_16440; // @[Mux.scala 19:72:@8446.4]
  wire [7:0] _T_16442; // @[Mux.scala 19:72:@8447.4]
  wire [7:0] _T_16449; // @[Mux.scala 19:72:@8454.4]
  wire [7:0] _T_16451; // @[Mux.scala 19:72:@8455.4]
  wire [7:0] _T_16452; // @[Mux.scala 19:72:@8456.4]
  wire [7:0] _T_16453; // @[Mux.scala 19:72:@8457.4]
  wire [7:0] _T_16454; // @[Mux.scala 19:72:@8458.4]
  wire [7:0] _T_16455; // @[Mux.scala 19:72:@8459.4]
  wire [7:0] _T_16456; // @[Mux.scala 19:72:@8460.4]
  wire [7:0] _T_16457; // @[Mux.scala 19:72:@8461.4]
  wire [7:0] _T_16458; // @[Mux.scala 19:72:@8462.4]
  wire [7:0] _T_16700; // @[Mux.scala 19:72:@8580.4]
  wire [7:0] _T_16702; // @[Mux.scala 19:72:@8581.4]
  wire [7:0] _T_16709; // @[Mux.scala 19:72:@8588.4]
  wire [7:0] _T_16711; // @[Mux.scala 19:72:@8589.4]
  wire [7:0] _T_16718; // @[Mux.scala 19:72:@8596.4]
  wire [7:0] _T_16720; // @[Mux.scala 19:72:@8597.4]
  wire [7:0] _T_16727; // @[Mux.scala 19:72:@8604.4]
  wire [7:0] _T_16729; // @[Mux.scala 19:72:@8605.4]
  wire [7:0] _T_16736; // @[Mux.scala 19:72:@8612.4]
  wire [7:0] _T_16738; // @[Mux.scala 19:72:@8613.4]
  wire [7:0] _T_16745; // @[Mux.scala 19:72:@8620.4]
  wire [7:0] _T_16747; // @[Mux.scala 19:72:@8621.4]
  wire [7:0] _T_16754; // @[Mux.scala 19:72:@8628.4]
  wire [7:0] _T_16756; // @[Mux.scala 19:72:@8629.4]
  wire [7:0] _T_16763; // @[Mux.scala 19:72:@8636.4]
  wire [7:0] _T_16765; // @[Mux.scala 19:72:@8637.4]
  wire [7:0] _T_16766; // @[Mux.scala 19:72:@8638.4]
  wire [7:0] _T_16767; // @[Mux.scala 19:72:@8639.4]
  wire [7:0] _T_16768; // @[Mux.scala 19:72:@8640.4]
  wire [7:0] _T_16769; // @[Mux.scala 19:72:@8641.4]
  wire [7:0] _T_16770; // @[Mux.scala 19:72:@8642.4]
  wire [7:0] _T_16771; // @[Mux.scala 19:72:@8643.4]
  wire [7:0] _T_16772; // @[Mux.scala 19:72:@8644.4]
  reg  storeAddrNotKnownFlagsPReg_0_0; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_147;
  reg  storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_148;
  reg  storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_149;
  reg  storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_150;
  reg  storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_151;
  reg  storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_152;
  reg  storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_153;
  reg  storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_154;
  reg  storeAddrNotKnownFlagsPReg_1_0; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_155;
  reg  storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_156;
  reg  storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_157;
  reg  storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_158;
  reg  storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_159;
  reg  storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_160;
  reg  storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_161;
  reg  storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_162;
  reg  storeAddrNotKnownFlagsPReg_2_0; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_163;
  reg  storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_164;
  reg  storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_165;
  reg  storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_166;
  reg  storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_167;
  reg  storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_168;
  reg  storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_169;
  reg  storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_170;
  reg  storeAddrNotKnownFlagsPReg_3_0; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_171;
  reg  storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_172;
  reg  storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_173;
  reg  storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_174;
  reg  storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_175;
  reg  storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_176;
  reg  storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_177;
  reg  storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_178;
  reg  storeAddrNotKnownFlagsPReg_4_0; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_179;
  reg  storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_180;
  reg  storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_181;
  reg  storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_182;
  reg  storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_183;
  reg  storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_184;
  reg  storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_185;
  reg  storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_186;
  reg  storeAddrNotKnownFlagsPReg_5_0; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_187;
  reg  storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_188;
  reg  storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_189;
  reg  storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_190;
  reg  storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_191;
  reg  storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_192;
  reg  storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_193;
  reg  storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_194;
  reg  storeAddrNotKnownFlagsPReg_6_0; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_195;
  reg  storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_196;
  reg  storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_197;
  reg  storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_198;
  reg  storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_199;
  reg  storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_200;
  reg  storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_201;
  reg  storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_202;
  reg  storeAddrNotKnownFlagsPReg_7_0; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_203;
  reg  storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_204;
  reg  storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_205;
  reg  storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_206;
  reg  storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_207;
  reg  storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_208;
  reg  storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_209;
  reg  storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 167:43:@8729.4]
  reg [31:0] _RAND_210;
  reg  shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 168:42:@8794.4]
  reg [31:0] _RAND_211;
  reg  shiftedStoreDataKnownPReg_1; // @[LoadQueue.scala 168:42:@8794.4]
  reg [31:0] _RAND_212;
  reg  shiftedStoreDataKnownPReg_2; // @[LoadQueue.scala 168:42:@8794.4]
  reg [31:0] _RAND_213;
  reg  shiftedStoreDataKnownPReg_3; // @[LoadQueue.scala 168:42:@8794.4]
  reg [31:0] _RAND_214;
  reg  shiftedStoreDataKnownPReg_4; // @[LoadQueue.scala 168:42:@8794.4]
  reg [31:0] _RAND_215;
  reg  shiftedStoreDataKnownPReg_5; // @[LoadQueue.scala 168:42:@8794.4]
  reg [31:0] _RAND_216;
  reg  shiftedStoreDataKnownPReg_6; // @[LoadQueue.scala 168:42:@8794.4]
  reg [31:0] _RAND_217;
  reg  shiftedStoreDataKnownPReg_7; // @[LoadQueue.scala 168:42:@8794.4]
  reg [31:0] _RAND_218;
  reg [31:0] shiftedStoreDataQPreg_0; // @[LoadQueue.scala 169:38:@8803.4]
  reg [31:0] _RAND_219;
  reg [31:0] shiftedStoreDataQPreg_1; // @[LoadQueue.scala 169:38:@8803.4]
  reg [31:0] _RAND_220;
  reg [31:0] shiftedStoreDataQPreg_2; // @[LoadQueue.scala 169:38:@8803.4]
  reg [31:0] _RAND_221;
  reg [31:0] shiftedStoreDataQPreg_3; // @[LoadQueue.scala 169:38:@8803.4]
  reg [31:0] _RAND_222;
  reg [31:0] shiftedStoreDataQPreg_4; // @[LoadQueue.scala 169:38:@8803.4]
  reg [31:0] _RAND_223;
  reg [31:0] shiftedStoreDataQPreg_5; // @[LoadQueue.scala 169:38:@8803.4]
  reg [31:0] _RAND_224;
  reg [31:0] shiftedStoreDataQPreg_6; // @[LoadQueue.scala 169:38:@8803.4]
  reg [31:0] _RAND_225;
  reg [31:0] shiftedStoreDataQPreg_7; // @[LoadQueue.scala 169:38:@8803.4]
  reg [31:0] _RAND_226;
  reg  addrKnownPReg_0; // @[LoadQueue.scala 170:30:@8812.4]
  reg [31:0] _RAND_227;
  reg  addrKnownPReg_1; // @[LoadQueue.scala 170:30:@8812.4]
  reg [31:0] _RAND_228;
  reg  addrKnownPReg_2; // @[LoadQueue.scala 170:30:@8812.4]
  reg [31:0] _RAND_229;
  reg  addrKnownPReg_3; // @[LoadQueue.scala 170:30:@8812.4]
  reg [31:0] _RAND_230;
  reg  addrKnownPReg_4; // @[LoadQueue.scala 170:30:@8812.4]
  reg [31:0] _RAND_231;
  reg  addrKnownPReg_5; // @[LoadQueue.scala 170:30:@8812.4]
  reg [31:0] _RAND_232;
  reg  addrKnownPReg_6; // @[LoadQueue.scala 170:30:@8812.4]
  reg [31:0] _RAND_233;
  reg  addrKnownPReg_7; // @[LoadQueue.scala 170:30:@8812.4]
  reg [31:0] _RAND_234;
  reg  dataKnownPReg_0; // @[LoadQueue.scala 171:30:@8821.4]
  reg [31:0] _RAND_235;
  reg  dataKnownPReg_1; // @[LoadQueue.scala 171:30:@8821.4]
  reg [31:0] _RAND_236;
  reg  dataKnownPReg_2; // @[LoadQueue.scala 171:30:@8821.4]
  reg [31:0] _RAND_237;
  reg  dataKnownPReg_3; // @[LoadQueue.scala 171:30:@8821.4]
  reg [31:0] _RAND_238;
  reg  dataKnownPReg_4; // @[LoadQueue.scala 171:30:@8821.4]
  reg [31:0] _RAND_239;
  reg  dataKnownPReg_5; // @[LoadQueue.scala 171:30:@8821.4]
  reg [31:0] _RAND_240;
  reg  dataKnownPReg_6; // @[LoadQueue.scala 171:30:@8821.4]
  reg [31:0] _RAND_241;
  reg  dataKnownPReg_7; // @[LoadQueue.scala 171:30:@8821.4]
  reg [31:0] _RAND_242;
  wire [1:0] _T_23532; // @[LoadQueue.scala 191:60:@8861.4]
  wire [1:0] _T_23533; // @[LoadQueue.scala 191:60:@8862.4]
  wire [2:0] _T_23534; // @[LoadQueue.scala 191:60:@8863.4]
  wire [2:0] _T_23535; // @[LoadQueue.scala 191:60:@8864.4]
  wire [2:0] _T_23536; // @[LoadQueue.scala 191:60:@8865.4]
  wire [2:0] _T_23537; // @[LoadQueue.scala 191:60:@8866.4]
  wire  _T_23540; // @[LoadQueue.scala 192:43:@8868.4]
  wire  _T_23541; // @[LoadQueue.scala 192:43:@8869.4]
  wire  _T_23542; // @[LoadQueue.scala 192:43:@8870.4]
  wire  _T_23543; // @[LoadQueue.scala 192:43:@8871.4]
  wire  _T_23544; // @[LoadQueue.scala 192:43:@8872.4]
  wire  _T_23545; // @[LoadQueue.scala 192:43:@8873.4]
  wire  _T_23546; // @[LoadQueue.scala 192:43:@8874.4]
  wire  _GEN_240; // @[LoadQueue.scala 193:43:@8876.6]
  wire  _GEN_241; // @[LoadQueue.scala 193:43:@8876.6]
  wire  _GEN_242; // @[LoadQueue.scala 193:43:@8876.6]
  wire  _GEN_243; // @[LoadQueue.scala 193:43:@8876.6]
  wire  _GEN_244; // @[LoadQueue.scala 193:43:@8876.6]
  wire  _GEN_245; // @[LoadQueue.scala 193:43:@8876.6]
  wire  _GEN_246; // @[LoadQueue.scala 193:43:@8876.6]
  wire  _GEN_247; // @[LoadQueue.scala 193:43:@8876.6]
  wire  _GEN_249; // @[LoadQueue.scala 194:31:@8877.6]
  wire  _GEN_250; // @[LoadQueue.scala 194:31:@8877.6]
  wire  _GEN_251; // @[LoadQueue.scala 194:31:@8877.6]
  wire  _GEN_252; // @[LoadQueue.scala 194:31:@8877.6]
  wire  _GEN_253; // @[LoadQueue.scala 194:31:@8877.6]
  wire  _GEN_254; // @[LoadQueue.scala 194:31:@8877.6]
  wire  _GEN_255; // @[LoadQueue.scala 194:31:@8877.6]
  wire [31:0] _GEN_257; // @[LoadQueue.scala 195:31:@8878.6]
  wire [31:0] _GEN_258; // @[LoadQueue.scala 195:31:@8878.6]
  wire [31:0] _GEN_259; // @[LoadQueue.scala 195:31:@8878.6]
  wire [31:0] _GEN_260; // @[LoadQueue.scala 195:31:@8878.6]
  wire [31:0] _GEN_261; // @[LoadQueue.scala 195:31:@8878.6]
  wire [31:0] _GEN_262; // @[LoadQueue.scala 195:31:@8878.6]
  wire [31:0] _GEN_263; // @[LoadQueue.scala 195:31:@8878.6]
  wire  lastConflict_0_0; // @[LoadQueue.scala 192:53:@8875.4]
  wire  lastConflict_0_1; // @[LoadQueue.scala 192:53:@8875.4]
  wire  lastConflict_0_2; // @[LoadQueue.scala 192:53:@8875.4]
  wire  lastConflict_0_3; // @[LoadQueue.scala 192:53:@8875.4]
  wire  lastConflict_0_4; // @[LoadQueue.scala 192:53:@8875.4]
  wire  lastConflict_0_5; // @[LoadQueue.scala 192:53:@8875.4]
  wire  lastConflict_0_6; // @[LoadQueue.scala 192:53:@8875.4]
  wire  lastConflict_0_7; // @[LoadQueue.scala 192:53:@8875.4]
  wire  canBypass_0; // @[LoadQueue.scala 192:53:@8875.4]
  wire [31:0] bypassVal_0; // @[LoadQueue.scala 192:53:@8875.4]
  wire [1:0] _T_23612; // @[LoadQueue.scala 191:60:@8908.4]
  wire [1:0] _T_23613; // @[LoadQueue.scala 191:60:@8909.4]
  wire [2:0] _T_23614; // @[LoadQueue.scala 191:60:@8910.4]
  wire [2:0] _T_23615; // @[LoadQueue.scala 191:60:@8911.4]
  wire [2:0] _T_23616; // @[LoadQueue.scala 191:60:@8912.4]
  wire [2:0] _T_23617; // @[LoadQueue.scala 191:60:@8913.4]
  wire  _T_23620; // @[LoadQueue.scala 192:43:@8915.4]
  wire  _T_23621; // @[LoadQueue.scala 192:43:@8916.4]
  wire  _T_23622; // @[LoadQueue.scala 192:43:@8917.4]
  wire  _T_23623; // @[LoadQueue.scala 192:43:@8918.4]
  wire  _T_23624; // @[LoadQueue.scala 192:43:@8919.4]
  wire  _T_23625; // @[LoadQueue.scala 192:43:@8920.4]
  wire  _T_23626; // @[LoadQueue.scala 192:43:@8921.4]
  wire  _GEN_274; // @[LoadQueue.scala 193:43:@8923.6]
  wire  _GEN_275; // @[LoadQueue.scala 193:43:@8923.6]
  wire  _GEN_276; // @[LoadQueue.scala 193:43:@8923.6]
  wire  _GEN_277; // @[LoadQueue.scala 193:43:@8923.6]
  wire  _GEN_278; // @[LoadQueue.scala 193:43:@8923.6]
  wire  _GEN_279; // @[LoadQueue.scala 193:43:@8923.6]
  wire  _GEN_280; // @[LoadQueue.scala 193:43:@8923.6]
  wire  _GEN_281; // @[LoadQueue.scala 193:43:@8923.6]
  wire  _GEN_283; // @[LoadQueue.scala 194:31:@8924.6]
  wire  _GEN_284; // @[LoadQueue.scala 194:31:@8924.6]
  wire  _GEN_285; // @[LoadQueue.scala 194:31:@8924.6]
  wire  _GEN_286; // @[LoadQueue.scala 194:31:@8924.6]
  wire  _GEN_287; // @[LoadQueue.scala 194:31:@8924.6]
  wire  _GEN_288; // @[LoadQueue.scala 194:31:@8924.6]
  wire  _GEN_289; // @[LoadQueue.scala 194:31:@8924.6]
  wire [31:0] _GEN_291; // @[LoadQueue.scala 195:31:@8925.6]
  wire [31:0] _GEN_292; // @[LoadQueue.scala 195:31:@8925.6]
  wire [31:0] _GEN_293; // @[LoadQueue.scala 195:31:@8925.6]
  wire [31:0] _GEN_294; // @[LoadQueue.scala 195:31:@8925.6]
  wire [31:0] _GEN_295; // @[LoadQueue.scala 195:31:@8925.6]
  wire [31:0] _GEN_296; // @[LoadQueue.scala 195:31:@8925.6]
  wire [31:0] _GEN_297; // @[LoadQueue.scala 195:31:@8925.6]
  wire  lastConflict_1_0; // @[LoadQueue.scala 192:53:@8922.4]
  wire  lastConflict_1_1; // @[LoadQueue.scala 192:53:@8922.4]
  wire  lastConflict_1_2; // @[LoadQueue.scala 192:53:@8922.4]
  wire  lastConflict_1_3; // @[LoadQueue.scala 192:53:@8922.4]
  wire  lastConflict_1_4; // @[LoadQueue.scala 192:53:@8922.4]
  wire  lastConflict_1_5; // @[LoadQueue.scala 192:53:@8922.4]
  wire  lastConflict_1_6; // @[LoadQueue.scala 192:53:@8922.4]
  wire  lastConflict_1_7; // @[LoadQueue.scala 192:53:@8922.4]
  wire  canBypass_1; // @[LoadQueue.scala 192:53:@8922.4]
  wire [31:0] bypassVal_1; // @[LoadQueue.scala 192:53:@8922.4]
  wire [1:0] _T_23692; // @[LoadQueue.scala 191:60:@8955.4]
  wire [1:0] _T_23693; // @[LoadQueue.scala 191:60:@8956.4]
  wire [2:0] _T_23694; // @[LoadQueue.scala 191:60:@8957.4]
  wire [2:0] _T_23695; // @[LoadQueue.scala 191:60:@8958.4]
  wire [2:0] _T_23696; // @[LoadQueue.scala 191:60:@8959.4]
  wire [2:0] _T_23697; // @[LoadQueue.scala 191:60:@8960.4]
  wire  _T_23700; // @[LoadQueue.scala 192:43:@8962.4]
  wire  _T_23701; // @[LoadQueue.scala 192:43:@8963.4]
  wire  _T_23702; // @[LoadQueue.scala 192:43:@8964.4]
  wire  _T_23703; // @[LoadQueue.scala 192:43:@8965.4]
  wire  _T_23704; // @[LoadQueue.scala 192:43:@8966.4]
  wire  _T_23705; // @[LoadQueue.scala 192:43:@8967.4]
  wire  _T_23706; // @[LoadQueue.scala 192:43:@8968.4]
  wire  _GEN_308; // @[LoadQueue.scala 193:43:@8970.6]
  wire  _GEN_309; // @[LoadQueue.scala 193:43:@8970.6]
  wire  _GEN_310; // @[LoadQueue.scala 193:43:@8970.6]
  wire  _GEN_311; // @[LoadQueue.scala 193:43:@8970.6]
  wire  _GEN_312; // @[LoadQueue.scala 193:43:@8970.6]
  wire  _GEN_313; // @[LoadQueue.scala 193:43:@8970.6]
  wire  _GEN_314; // @[LoadQueue.scala 193:43:@8970.6]
  wire  _GEN_315; // @[LoadQueue.scala 193:43:@8970.6]
  wire  _GEN_317; // @[LoadQueue.scala 194:31:@8971.6]
  wire  _GEN_318; // @[LoadQueue.scala 194:31:@8971.6]
  wire  _GEN_319; // @[LoadQueue.scala 194:31:@8971.6]
  wire  _GEN_320; // @[LoadQueue.scala 194:31:@8971.6]
  wire  _GEN_321; // @[LoadQueue.scala 194:31:@8971.6]
  wire  _GEN_322; // @[LoadQueue.scala 194:31:@8971.6]
  wire  _GEN_323; // @[LoadQueue.scala 194:31:@8971.6]
  wire [31:0] _GEN_325; // @[LoadQueue.scala 195:31:@8972.6]
  wire [31:0] _GEN_326; // @[LoadQueue.scala 195:31:@8972.6]
  wire [31:0] _GEN_327; // @[LoadQueue.scala 195:31:@8972.6]
  wire [31:0] _GEN_328; // @[LoadQueue.scala 195:31:@8972.6]
  wire [31:0] _GEN_329; // @[LoadQueue.scala 195:31:@8972.6]
  wire [31:0] _GEN_330; // @[LoadQueue.scala 195:31:@8972.6]
  wire [31:0] _GEN_331; // @[LoadQueue.scala 195:31:@8972.6]
  wire  lastConflict_2_0; // @[LoadQueue.scala 192:53:@8969.4]
  wire  lastConflict_2_1; // @[LoadQueue.scala 192:53:@8969.4]
  wire  lastConflict_2_2; // @[LoadQueue.scala 192:53:@8969.4]
  wire  lastConflict_2_3; // @[LoadQueue.scala 192:53:@8969.4]
  wire  lastConflict_2_4; // @[LoadQueue.scala 192:53:@8969.4]
  wire  lastConflict_2_5; // @[LoadQueue.scala 192:53:@8969.4]
  wire  lastConflict_2_6; // @[LoadQueue.scala 192:53:@8969.4]
  wire  lastConflict_2_7; // @[LoadQueue.scala 192:53:@8969.4]
  wire  canBypass_2; // @[LoadQueue.scala 192:53:@8969.4]
  wire [31:0] bypassVal_2; // @[LoadQueue.scala 192:53:@8969.4]
  wire [1:0] _T_23772; // @[LoadQueue.scala 191:60:@9002.4]
  wire [1:0] _T_23773; // @[LoadQueue.scala 191:60:@9003.4]
  wire [2:0] _T_23774; // @[LoadQueue.scala 191:60:@9004.4]
  wire [2:0] _T_23775; // @[LoadQueue.scala 191:60:@9005.4]
  wire [2:0] _T_23776; // @[LoadQueue.scala 191:60:@9006.4]
  wire [2:0] _T_23777; // @[LoadQueue.scala 191:60:@9007.4]
  wire  _T_23780; // @[LoadQueue.scala 192:43:@9009.4]
  wire  _T_23781; // @[LoadQueue.scala 192:43:@9010.4]
  wire  _T_23782; // @[LoadQueue.scala 192:43:@9011.4]
  wire  _T_23783; // @[LoadQueue.scala 192:43:@9012.4]
  wire  _T_23784; // @[LoadQueue.scala 192:43:@9013.4]
  wire  _T_23785; // @[LoadQueue.scala 192:43:@9014.4]
  wire  _T_23786; // @[LoadQueue.scala 192:43:@9015.4]
  wire  _GEN_342; // @[LoadQueue.scala 193:43:@9017.6]
  wire  _GEN_343; // @[LoadQueue.scala 193:43:@9017.6]
  wire  _GEN_344; // @[LoadQueue.scala 193:43:@9017.6]
  wire  _GEN_345; // @[LoadQueue.scala 193:43:@9017.6]
  wire  _GEN_346; // @[LoadQueue.scala 193:43:@9017.6]
  wire  _GEN_347; // @[LoadQueue.scala 193:43:@9017.6]
  wire  _GEN_348; // @[LoadQueue.scala 193:43:@9017.6]
  wire  _GEN_349; // @[LoadQueue.scala 193:43:@9017.6]
  wire  _GEN_351; // @[LoadQueue.scala 194:31:@9018.6]
  wire  _GEN_352; // @[LoadQueue.scala 194:31:@9018.6]
  wire  _GEN_353; // @[LoadQueue.scala 194:31:@9018.6]
  wire  _GEN_354; // @[LoadQueue.scala 194:31:@9018.6]
  wire  _GEN_355; // @[LoadQueue.scala 194:31:@9018.6]
  wire  _GEN_356; // @[LoadQueue.scala 194:31:@9018.6]
  wire  _GEN_357; // @[LoadQueue.scala 194:31:@9018.6]
  wire [31:0] _GEN_359; // @[LoadQueue.scala 195:31:@9019.6]
  wire [31:0] _GEN_360; // @[LoadQueue.scala 195:31:@9019.6]
  wire [31:0] _GEN_361; // @[LoadQueue.scala 195:31:@9019.6]
  wire [31:0] _GEN_362; // @[LoadQueue.scala 195:31:@9019.6]
  wire [31:0] _GEN_363; // @[LoadQueue.scala 195:31:@9019.6]
  wire [31:0] _GEN_364; // @[LoadQueue.scala 195:31:@9019.6]
  wire [31:0] _GEN_365; // @[LoadQueue.scala 195:31:@9019.6]
  wire  lastConflict_3_0; // @[LoadQueue.scala 192:53:@9016.4]
  wire  lastConflict_3_1; // @[LoadQueue.scala 192:53:@9016.4]
  wire  lastConflict_3_2; // @[LoadQueue.scala 192:53:@9016.4]
  wire  lastConflict_3_3; // @[LoadQueue.scala 192:53:@9016.4]
  wire  lastConflict_3_4; // @[LoadQueue.scala 192:53:@9016.4]
  wire  lastConflict_3_5; // @[LoadQueue.scala 192:53:@9016.4]
  wire  lastConflict_3_6; // @[LoadQueue.scala 192:53:@9016.4]
  wire  lastConflict_3_7; // @[LoadQueue.scala 192:53:@9016.4]
  wire  canBypass_3; // @[LoadQueue.scala 192:53:@9016.4]
  wire [31:0] bypassVal_3; // @[LoadQueue.scala 192:53:@9016.4]
  wire [1:0] _T_23852; // @[LoadQueue.scala 191:60:@9049.4]
  wire [1:0] _T_23853; // @[LoadQueue.scala 191:60:@9050.4]
  wire [2:0] _T_23854; // @[LoadQueue.scala 191:60:@9051.4]
  wire [2:0] _T_23855; // @[LoadQueue.scala 191:60:@9052.4]
  wire [2:0] _T_23856; // @[LoadQueue.scala 191:60:@9053.4]
  wire [2:0] _T_23857; // @[LoadQueue.scala 191:60:@9054.4]
  wire  _T_23860; // @[LoadQueue.scala 192:43:@9056.4]
  wire  _T_23861; // @[LoadQueue.scala 192:43:@9057.4]
  wire  _T_23862; // @[LoadQueue.scala 192:43:@9058.4]
  wire  _T_23863; // @[LoadQueue.scala 192:43:@9059.4]
  wire  _T_23864; // @[LoadQueue.scala 192:43:@9060.4]
  wire  _T_23865; // @[LoadQueue.scala 192:43:@9061.4]
  wire  _T_23866; // @[LoadQueue.scala 192:43:@9062.4]
  wire  _GEN_376; // @[LoadQueue.scala 193:43:@9064.6]
  wire  _GEN_377; // @[LoadQueue.scala 193:43:@9064.6]
  wire  _GEN_378; // @[LoadQueue.scala 193:43:@9064.6]
  wire  _GEN_379; // @[LoadQueue.scala 193:43:@9064.6]
  wire  _GEN_380; // @[LoadQueue.scala 193:43:@9064.6]
  wire  _GEN_381; // @[LoadQueue.scala 193:43:@9064.6]
  wire  _GEN_382; // @[LoadQueue.scala 193:43:@9064.6]
  wire  _GEN_383; // @[LoadQueue.scala 193:43:@9064.6]
  wire  _GEN_385; // @[LoadQueue.scala 194:31:@9065.6]
  wire  _GEN_386; // @[LoadQueue.scala 194:31:@9065.6]
  wire  _GEN_387; // @[LoadQueue.scala 194:31:@9065.6]
  wire  _GEN_388; // @[LoadQueue.scala 194:31:@9065.6]
  wire  _GEN_389; // @[LoadQueue.scala 194:31:@9065.6]
  wire  _GEN_390; // @[LoadQueue.scala 194:31:@9065.6]
  wire  _GEN_391; // @[LoadQueue.scala 194:31:@9065.6]
  wire [31:0] _GEN_393; // @[LoadQueue.scala 195:31:@9066.6]
  wire [31:0] _GEN_394; // @[LoadQueue.scala 195:31:@9066.6]
  wire [31:0] _GEN_395; // @[LoadQueue.scala 195:31:@9066.6]
  wire [31:0] _GEN_396; // @[LoadQueue.scala 195:31:@9066.6]
  wire [31:0] _GEN_397; // @[LoadQueue.scala 195:31:@9066.6]
  wire [31:0] _GEN_398; // @[LoadQueue.scala 195:31:@9066.6]
  wire [31:0] _GEN_399; // @[LoadQueue.scala 195:31:@9066.6]
  wire  lastConflict_4_0; // @[LoadQueue.scala 192:53:@9063.4]
  wire  lastConflict_4_1; // @[LoadQueue.scala 192:53:@9063.4]
  wire  lastConflict_4_2; // @[LoadQueue.scala 192:53:@9063.4]
  wire  lastConflict_4_3; // @[LoadQueue.scala 192:53:@9063.4]
  wire  lastConflict_4_4; // @[LoadQueue.scala 192:53:@9063.4]
  wire  lastConflict_4_5; // @[LoadQueue.scala 192:53:@9063.4]
  wire  lastConflict_4_6; // @[LoadQueue.scala 192:53:@9063.4]
  wire  lastConflict_4_7; // @[LoadQueue.scala 192:53:@9063.4]
  wire  canBypass_4; // @[LoadQueue.scala 192:53:@9063.4]
  wire [31:0] bypassVal_4; // @[LoadQueue.scala 192:53:@9063.4]
  wire [1:0] _T_23932; // @[LoadQueue.scala 191:60:@9096.4]
  wire [1:0] _T_23933; // @[LoadQueue.scala 191:60:@9097.4]
  wire [2:0] _T_23934; // @[LoadQueue.scala 191:60:@9098.4]
  wire [2:0] _T_23935; // @[LoadQueue.scala 191:60:@9099.4]
  wire [2:0] _T_23936; // @[LoadQueue.scala 191:60:@9100.4]
  wire [2:0] _T_23937; // @[LoadQueue.scala 191:60:@9101.4]
  wire  _T_23940; // @[LoadQueue.scala 192:43:@9103.4]
  wire  _T_23941; // @[LoadQueue.scala 192:43:@9104.4]
  wire  _T_23942; // @[LoadQueue.scala 192:43:@9105.4]
  wire  _T_23943; // @[LoadQueue.scala 192:43:@9106.4]
  wire  _T_23944; // @[LoadQueue.scala 192:43:@9107.4]
  wire  _T_23945; // @[LoadQueue.scala 192:43:@9108.4]
  wire  _T_23946; // @[LoadQueue.scala 192:43:@9109.4]
  wire  _GEN_410; // @[LoadQueue.scala 193:43:@9111.6]
  wire  _GEN_411; // @[LoadQueue.scala 193:43:@9111.6]
  wire  _GEN_412; // @[LoadQueue.scala 193:43:@9111.6]
  wire  _GEN_413; // @[LoadQueue.scala 193:43:@9111.6]
  wire  _GEN_414; // @[LoadQueue.scala 193:43:@9111.6]
  wire  _GEN_415; // @[LoadQueue.scala 193:43:@9111.6]
  wire  _GEN_416; // @[LoadQueue.scala 193:43:@9111.6]
  wire  _GEN_417; // @[LoadQueue.scala 193:43:@9111.6]
  wire  _GEN_419; // @[LoadQueue.scala 194:31:@9112.6]
  wire  _GEN_420; // @[LoadQueue.scala 194:31:@9112.6]
  wire  _GEN_421; // @[LoadQueue.scala 194:31:@9112.6]
  wire  _GEN_422; // @[LoadQueue.scala 194:31:@9112.6]
  wire  _GEN_423; // @[LoadQueue.scala 194:31:@9112.6]
  wire  _GEN_424; // @[LoadQueue.scala 194:31:@9112.6]
  wire  _GEN_425; // @[LoadQueue.scala 194:31:@9112.6]
  wire [31:0] _GEN_427; // @[LoadQueue.scala 195:31:@9113.6]
  wire [31:0] _GEN_428; // @[LoadQueue.scala 195:31:@9113.6]
  wire [31:0] _GEN_429; // @[LoadQueue.scala 195:31:@9113.6]
  wire [31:0] _GEN_430; // @[LoadQueue.scala 195:31:@9113.6]
  wire [31:0] _GEN_431; // @[LoadQueue.scala 195:31:@9113.6]
  wire [31:0] _GEN_432; // @[LoadQueue.scala 195:31:@9113.6]
  wire [31:0] _GEN_433; // @[LoadQueue.scala 195:31:@9113.6]
  wire  lastConflict_5_0; // @[LoadQueue.scala 192:53:@9110.4]
  wire  lastConflict_5_1; // @[LoadQueue.scala 192:53:@9110.4]
  wire  lastConflict_5_2; // @[LoadQueue.scala 192:53:@9110.4]
  wire  lastConflict_5_3; // @[LoadQueue.scala 192:53:@9110.4]
  wire  lastConflict_5_4; // @[LoadQueue.scala 192:53:@9110.4]
  wire  lastConflict_5_5; // @[LoadQueue.scala 192:53:@9110.4]
  wire  lastConflict_5_6; // @[LoadQueue.scala 192:53:@9110.4]
  wire  lastConflict_5_7; // @[LoadQueue.scala 192:53:@9110.4]
  wire  canBypass_5; // @[LoadQueue.scala 192:53:@9110.4]
  wire [31:0] bypassVal_5; // @[LoadQueue.scala 192:53:@9110.4]
  wire [1:0] _T_24012; // @[LoadQueue.scala 191:60:@9143.4]
  wire [1:0] _T_24013; // @[LoadQueue.scala 191:60:@9144.4]
  wire [2:0] _T_24014; // @[LoadQueue.scala 191:60:@9145.4]
  wire [2:0] _T_24015; // @[LoadQueue.scala 191:60:@9146.4]
  wire [2:0] _T_24016; // @[LoadQueue.scala 191:60:@9147.4]
  wire [2:0] _T_24017; // @[LoadQueue.scala 191:60:@9148.4]
  wire  _T_24020; // @[LoadQueue.scala 192:43:@9150.4]
  wire  _T_24021; // @[LoadQueue.scala 192:43:@9151.4]
  wire  _T_24022; // @[LoadQueue.scala 192:43:@9152.4]
  wire  _T_24023; // @[LoadQueue.scala 192:43:@9153.4]
  wire  _T_24024; // @[LoadQueue.scala 192:43:@9154.4]
  wire  _T_24025; // @[LoadQueue.scala 192:43:@9155.4]
  wire  _T_24026; // @[LoadQueue.scala 192:43:@9156.4]
  wire  _GEN_444; // @[LoadQueue.scala 193:43:@9158.6]
  wire  _GEN_445; // @[LoadQueue.scala 193:43:@9158.6]
  wire  _GEN_446; // @[LoadQueue.scala 193:43:@9158.6]
  wire  _GEN_447; // @[LoadQueue.scala 193:43:@9158.6]
  wire  _GEN_448; // @[LoadQueue.scala 193:43:@9158.6]
  wire  _GEN_449; // @[LoadQueue.scala 193:43:@9158.6]
  wire  _GEN_450; // @[LoadQueue.scala 193:43:@9158.6]
  wire  _GEN_451; // @[LoadQueue.scala 193:43:@9158.6]
  wire  _GEN_453; // @[LoadQueue.scala 194:31:@9159.6]
  wire  _GEN_454; // @[LoadQueue.scala 194:31:@9159.6]
  wire  _GEN_455; // @[LoadQueue.scala 194:31:@9159.6]
  wire  _GEN_456; // @[LoadQueue.scala 194:31:@9159.6]
  wire  _GEN_457; // @[LoadQueue.scala 194:31:@9159.6]
  wire  _GEN_458; // @[LoadQueue.scala 194:31:@9159.6]
  wire  _GEN_459; // @[LoadQueue.scala 194:31:@9159.6]
  wire [31:0] _GEN_461; // @[LoadQueue.scala 195:31:@9160.6]
  wire [31:0] _GEN_462; // @[LoadQueue.scala 195:31:@9160.6]
  wire [31:0] _GEN_463; // @[LoadQueue.scala 195:31:@9160.6]
  wire [31:0] _GEN_464; // @[LoadQueue.scala 195:31:@9160.6]
  wire [31:0] _GEN_465; // @[LoadQueue.scala 195:31:@9160.6]
  wire [31:0] _GEN_466; // @[LoadQueue.scala 195:31:@9160.6]
  wire [31:0] _GEN_467; // @[LoadQueue.scala 195:31:@9160.6]
  wire  lastConflict_6_0; // @[LoadQueue.scala 192:53:@9157.4]
  wire  lastConflict_6_1; // @[LoadQueue.scala 192:53:@9157.4]
  wire  lastConflict_6_2; // @[LoadQueue.scala 192:53:@9157.4]
  wire  lastConflict_6_3; // @[LoadQueue.scala 192:53:@9157.4]
  wire  lastConflict_6_4; // @[LoadQueue.scala 192:53:@9157.4]
  wire  lastConflict_6_5; // @[LoadQueue.scala 192:53:@9157.4]
  wire  lastConflict_6_6; // @[LoadQueue.scala 192:53:@9157.4]
  wire  lastConflict_6_7; // @[LoadQueue.scala 192:53:@9157.4]
  wire  canBypass_6; // @[LoadQueue.scala 192:53:@9157.4]
  wire [31:0] bypassVal_6; // @[LoadQueue.scala 192:53:@9157.4]
  wire [1:0] _T_24092; // @[LoadQueue.scala 191:60:@9190.4]
  wire [1:0] _T_24093; // @[LoadQueue.scala 191:60:@9191.4]
  wire [2:0] _T_24094; // @[LoadQueue.scala 191:60:@9192.4]
  wire [2:0] _T_24095; // @[LoadQueue.scala 191:60:@9193.4]
  wire [2:0] _T_24096; // @[LoadQueue.scala 191:60:@9194.4]
  wire [2:0] _T_24097; // @[LoadQueue.scala 191:60:@9195.4]
  wire  _T_24100; // @[LoadQueue.scala 192:43:@9197.4]
  wire  _T_24101; // @[LoadQueue.scala 192:43:@9198.4]
  wire  _T_24102; // @[LoadQueue.scala 192:43:@9199.4]
  wire  _T_24103; // @[LoadQueue.scala 192:43:@9200.4]
  wire  _T_24104; // @[LoadQueue.scala 192:43:@9201.4]
  wire  _T_24105; // @[LoadQueue.scala 192:43:@9202.4]
  wire  _T_24106; // @[LoadQueue.scala 192:43:@9203.4]
  wire  _GEN_478; // @[LoadQueue.scala 193:43:@9205.6]
  wire  _GEN_479; // @[LoadQueue.scala 193:43:@9205.6]
  wire  _GEN_480; // @[LoadQueue.scala 193:43:@9205.6]
  wire  _GEN_481; // @[LoadQueue.scala 193:43:@9205.6]
  wire  _GEN_482; // @[LoadQueue.scala 193:43:@9205.6]
  wire  _GEN_483; // @[LoadQueue.scala 193:43:@9205.6]
  wire  _GEN_484; // @[LoadQueue.scala 193:43:@9205.6]
  wire  _GEN_485; // @[LoadQueue.scala 193:43:@9205.6]
  wire  _GEN_487; // @[LoadQueue.scala 194:31:@9206.6]
  wire  _GEN_488; // @[LoadQueue.scala 194:31:@9206.6]
  wire  _GEN_489; // @[LoadQueue.scala 194:31:@9206.6]
  wire  _GEN_490; // @[LoadQueue.scala 194:31:@9206.6]
  wire  _GEN_491; // @[LoadQueue.scala 194:31:@9206.6]
  wire  _GEN_492; // @[LoadQueue.scala 194:31:@9206.6]
  wire  _GEN_493; // @[LoadQueue.scala 194:31:@9206.6]
  wire [31:0] _GEN_495; // @[LoadQueue.scala 195:31:@9207.6]
  wire [31:0] _GEN_496; // @[LoadQueue.scala 195:31:@9207.6]
  wire [31:0] _GEN_497; // @[LoadQueue.scala 195:31:@9207.6]
  wire [31:0] _GEN_498; // @[LoadQueue.scala 195:31:@9207.6]
  wire [31:0] _GEN_499; // @[LoadQueue.scala 195:31:@9207.6]
  wire [31:0] _GEN_500; // @[LoadQueue.scala 195:31:@9207.6]
  wire [31:0] _GEN_501; // @[LoadQueue.scala 195:31:@9207.6]
  wire  lastConflict_7_0; // @[LoadQueue.scala 192:53:@9204.4]
  wire  lastConflict_7_1; // @[LoadQueue.scala 192:53:@9204.4]
  wire  lastConflict_7_2; // @[LoadQueue.scala 192:53:@9204.4]
  wire  lastConflict_7_3; // @[LoadQueue.scala 192:53:@9204.4]
  wire  lastConflict_7_4; // @[LoadQueue.scala 192:53:@9204.4]
  wire  lastConflict_7_5; // @[LoadQueue.scala 192:53:@9204.4]
  wire  lastConflict_7_6; // @[LoadQueue.scala 192:53:@9204.4]
  wire  lastConflict_7_7; // @[LoadQueue.scala 192:53:@9204.4]
  wire  canBypass_7; // @[LoadQueue.scala 192:53:@9204.4]
  wire [31:0] bypassVal_7; // @[LoadQueue.scala 192:53:@9204.4]
  wire [7:0] _T_24150; // @[OneHot.scala 52:12:@9212.4]
  wire  _T_24152; // @[util.scala 33:60:@9214.4]
  wire  _T_24153; // @[util.scala 33:60:@9215.4]
  wire  _T_24154; // @[util.scala 33:60:@9216.4]
  wire  _T_24155; // @[util.scala 33:60:@9217.4]
  wire  _T_24156; // @[util.scala 33:60:@9218.4]
  wire  _T_24157; // @[util.scala 33:60:@9219.4]
  wire  _T_24158; // @[util.scala 33:60:@9220.4]
  wire  _T_24159; // @[util.scala 33:60:@9221.4]
  wire  _T_25144; // @[LoadQueue.scala 229:41:@9968.4]
  wire  _T_25145; // @[LoadQueue.scala 229:38:@9969.4]
  wire  _T_25147; // @[LoadQueue.scala 230:12:@9971.6]
  reg  prevPriorityRequest_7; // @[LoadQueue.scala 207:36:@9530.4]
  reg [31:0] _RAND_243;
  wire  _T_25149; // @[LoadQueue.scala 230:46:@9972.6]
  wire  _T_25150; // @[LoadQueue.scala 230:43:@9973.6]
  wire  _T_25152; // @[LoadQueue.scala 230:84:@9974.6]
  wire  _T_25153; // @[LoadQueue.scala 230:81:@9975.6]
  wire  _T_25156; // @[LoadQueue.scala 233:86:@9978.8]
  wire  _T_25157; // @[LoadQueue.scala 233:86:@9979.8]
  wire  _T_25158; // @[LoadQueue.scala 233:86:@9980.8]
  wire  _T_25159; // @[LoadQueue.scala 233:86:@9981.8]
  wire  _T_25160; // @[LoadQueue.scala 233:86:@9982.8]
  wire  _T_25161; // @[LoadQueue.scala 233:86:@9983.8]
  wire  _T_25162; // @[LoadQueue.scala 233:86:@9984.8]
  wire  _T_25164; // @[LoadQueue.scala 233:38:@9985.8]
  wire  _T_25175; // @[LoadQueue.scala 234:11:@9994.8]
  wire  _T_25176; // @[LoadQueue.scala 233:103:@9995.8]
  wire  _GEN_564; // @[LoadQueue.scala 230:110:@9976.6]
  wire  loadRequest_7; // @[LoadQueue.scala 229:71:@9970.4]
  wire [7:0] _T_24184; // @[Mux.scala 31:69:@9231.4]
  wire  _T_25092; // @[LoadQueue.scala 229:41:@9918.4]
  wire  _T_25093; // @[LoadQueue.scala 229:38:@9919.4]
  wire  _T_25095; // @[LoadQueue.scala 230:12:@9921.6]
  reg  prevPriorityRequest_6; // @[LoadQueue.scala 207:36:@9530.4]
  reg [31:0] _RAND_244;
  wire  _T_25097; // @[LoadQueue.scala 230:46:@9922.6]
  wire  _T_25098; // @[LoadQueue.scala 230:43:@9923.6]
  wire  _T_25100; // @[LoadQueue.scala 230:84:@9924.6]
  wire  _T_25101; // @[LoadQueue.scala 230:81:@9925.6]
  wire  _T_25104; // @[LoadQueue.scala 233:86:@9928.8]
  wire  _T_25105; // @[LoadQueue.scala 233:86:@9929.8]
  wire  _T_25106; // @[LoadQueue.scala 233:86:@9930.8]
  wire  _T_25107; // @[LoadQueue.scala 233:86:@9931.8]
  wire  _T_25108; // @[LoadQueue.scala 233:86:@9932.8]
  wire  _T_25109; // @[LoadQueue.scala 233:86:@9933.8]
  wire  _T_25110; // @[LoadQueue.scala 233:86:@9934.8]
  wire  _T_25112; // @[LoadQueue.scala 233:38:@9935.8]
  wire  _T_25123; // @[LoadQueue.scala 234:11:@9944.8]
  wire  _T_25124; // @[LoadQueue.scala 233:103:@9945.8]
  wire  _GEN_560; // @[LoadQueue.scala 230:110:@9926.6]
  wire  loadRequest_6; // @[LoadQueue.scala 229:71:@9920.4]
  wire [7:0] _T_24185; // @[Mux.scala 31:69:@9232.4]
  wire  _T_25040; // @[LoadQueue.scala 229:41:@9868.4]
  wire  _T_25041; // @[LoadQueue.scala 229:38:@9869.4]
  wire  _T_25043; // @[LoadQueue.scala 230:12:@9871.6]
  reg  prevPriorityRequest_5; // @[LoadQueue.scala 207:36:@9530.4]
  reg [31:0] _RAND_245;
  wire  _T_25045; // @[LoadQueue.scala 230:46:@9872.6]
  wire  _T_25046; // @[LoadQueue.scala 230:43:@9873.6]
  wire  _T_25048; // @[LoadQueue.scala 230:84:@9874.6]
  wire  _T_25049; // @[LoadQueue.scala 230:81:@9875.6]
  wire  _T_25052; // @[LoadQueue.scala 233:86:@9878.8]
  wire  _T_25053; // @[LoadQueue.scala 233:86:@9879.8]
  wire  _T_25054; // @[LoadQueue.scala 233:86:@9880.8]
  wire  _T_25055; // @[LoadQueue.scala 233:86:@9881.8]
  wire  _T_25056; // @[LoadQueue.scala 233:86:@9882.8]
  wire  _T_25057; // @[LoadQueue.scala 233:86:@9883.8]
  wire  _T_25058; // @[LoadQueue.scala 233:86:@9884.8]
  wire  _T_25060; // @[LoadQueue.scala 233:38:@9885.8]
  wire  _T_25071; // @[LoadQueue.scala 234:11:@9894.8]
  wire  _T_25072; // @[LoadQueue.scala 233:103:@9895.8]
  wire  _GEN_556; // @[LoadQueue.scala 230:110:@9876.6]
  wire  loadRequest_5; // @[LoadQueue.scala 229:71:@9870.4]
  wire [7:0] _T_24186; // @[Mux.scala 31:69:@9233.4]
  wire  _T_24988; // @[LoadQueue.scala 229:41:@9818.4]
  wire  _T_24989; // @[LoadQueue.scala 229:38:@9819.4]
  wire  _T_24991; // @[LoadQueue.scala 230:12:@9821.6]
  reg  prevPriorityRequest_4; // @[LoadQueue.scala 207:36:@9530.4]
  reg [31:0] _RAND_246;
  wire  _T_24993; // @[LoadQueue.scala 230:46:@9822.6]
  wire  _T_24994; // @[LoadQueue.scala 230:43:@9823.6]
  wire  _T_24996; // @[LoadQueue.scala 230:84:@9824.6]
  wire  _T_24997; // @[LoadQueue.scala 230:81:@9825.6]
  wire  _T_25000; // @[LoadQueue.scala 233:86:@9828.8]
  wire  _T_25001; // @[LoadQueue.scala 233:86:@9829.8]
  wire  _T_25002; // @[LoadQueue.scala 233:86:@9830.8]
  wire  _T_25003; // @[LoadQueue.scala 233:86:@9831.8]
  wire  _T_25004; // @[LoadQueue.scala 233:86:@9832.8]
  wire  _T_25005; // @[LoadQueue.scala 233:86:@9833.8]
  wire  _T_25006; // @[LoadQueue.scala 233:86:@9834.8]
  wire  _T_25008; // @[LoadQueue.scala 233:38:@9835.8]
  wire  _T_25019; // @[LoadQueue.scala 234:11:@9844.8]
  wire  _T_25020; // @[LoadQueue.scala 233:103:@9845.8]
  wire  _GEN_552; // @[LoadQueue.scala 230:110:@9826.6]
  wire  loadRequest_4; // @[LoadQueue.scala 229:71:@9820.4]
  wire [7:0] _T_24187; // @[Mux.scala 31:69:@9234.4]
  wire  _T_24936; // @[LoadQueue.scala 229:41:@9768.4]
  wire  _T_24937; // @[LoadQueue.scala 229:38:@9769.4]
  wire  _T_24939; // @[LoadQueue.scala 230:12:@9771.6]
  reg  prevPriorityRequest_3; // @[LoadQueue.scala 207:36:@9530.4]
  reg [31:0] _RAND_247;
  wire  _T_24941; // @[LoadQueue.scala 230:46:@9772.6]
  wire  _T_24942; // @[LoadQueue.scala 230:43:@9773.6]
  wire  _T_24944; // @[LoadQueue.scala 230:84:@9774.6]
  wire  _T_24945; // @[LoadQueue.scala 230:81:@9775.6]
  wire  _T_24948; // @[LoadQueue.scala 233:86:@9778.8]
  wire  _T_24949; // @[LoadQueue.scala 233:86:@9779.8]
  wire  _T_24950; // @[LoadQueue.scala 233:86:@9780.8]
  wire  _T_24951; // @[LoadQueue.scala 233:86:@9781.8]
  wire  _T_24952; // @[LoadQueue.scala 233:86:@9782.8]
  wire  _T_24953; // @[LoadQueue.scala 233:86:@9783.8]
  wire  _T_24954; // @[LoadQueue.scala 233:86:@9784.8]
  wire  _T_24956; // @[LoadQueue.scala 233:38:@9785.8]
  wire  _T_24967; // @[LoadQueue.scala 234:11:@9794.8]
  wire  _T_24968; // @[LoadQueue.scala 233:103:@9795.8]
  wire  _GEN_548; // @[LoadQueue.scala 230:110:@9776.6]
  wire  loadRequest_3; // @[LoadQueue.scala 229:71:@9770.4]
  wire [7:0] _T_24188; // @[Mux.scala 31:69:@9235.4]
  wire  _T_24884; // @[LoadQueue.scala 229:41:@9718.4]
  wire  _T_24885; // @[LoadQueue.scala 229:38:@9719.4]
  wire  _T_24887; // @[LoadQueue.scala 230:12:@9721.6]
  reg  prevPriorityRequest_2; // @[LoadQueue.scala 207:36:@9530.4]
  reg [31:0] _RAND_248;
  wire  _T_24889; // @[LoadQueue.scala 230:46:@9722.6]
  wire  _T_24890; // @[LoadQueue.scala 230:43:@9723.6]
  wire  _T_24892; // @[LoadQueue.scala 230:84:@9724.6]
  wire  _T_24893; // @[LoadQueue.scala 230:81:@9725.6]
  wire  _T_24896; // @[LoadQueue.scala 233:86:@9728.8]
  wire  _T_24897; // @[LoadQueue.scala 233:86:@9729.8]
  wire  _T_24898; // @[LoadQueue.scala 233:86:@9730.8]
  wire  _T_24899; // @[LoadQueue.scala 233:86:@9731.8]
  wire  _T_24900; // @[LoadQueue.scala 233:86:@9732.8]
  wire  _T_24901; // @[LoadQueue.scala 233:86:@9733.8]
  wire  _T_24902; // @[LoadQueue.scala 233:86:@9734.8]
  wire  _T_24904; // @[LoadQueue.scala 233:38:@9735.8]
  wire  _T_24915; // @[LoadQueue.scala 234:11:@9744.8]
  wire  _T_24916; // @[LoadQueue.scala 233:103:@9745.8]
  wire  _GEN_544; // @[LoadQueue.scala 230:110:@9726.6]
  wire  loadRequest_2; // @[LoadQueue.scala 229:71:@9720.4]
  wire [7:0] _T_24189; // @[Mux.scala 31:69:@9236.4]
  wire  _T_24832; // @[LoadQueue.scala 229:41:@9668.4]
  wire  _T_24833; // @[LoadQueue.scala 229:38:@9669.4]
  wire  _T_24835; // @[LoadQueue.scala 230:12:@9671.6]
  reg  prevPriorityRequest_1; // @[LoadQueue.scala 207:36:@9530.4]
  reg [31:0] _RAND_249;
  wire  _T_24837; // @[LoadQueue.scala 230:46:@9672.6]
  wire  _T_24838; // @[LoadQueue.scala 230:43:@9673.6]
  wire  _T_24840; // @[LoadQueue.scala 230:84:@9674.6]
  wire  _T_24841; // @[LoadQueue.scala 230:81:@9675.6]
  wire  _T_24844; // @[LoadQueue.scala 233:86:@9678.8]
  wire  _T_24845; // @[LoadQueue.scala 233:86:@9679.8]
  wire  _T_24846; // @[LoadQueue.scala 233:86:@9680.8]
  wire  _T_24847; // @[LoadQueue.scala 233:86:@9681.8]
  wire  _T_24848; // @[LoadQueue.scala 233:86:@9682.8]
  wire  _T_24849; // @[LoadQueue.scala 233:86:@9683.8]
  wire  _T_24850; // @[LoadQueue.scala 233:86:@9684.8]
  wire  _T_24852; // @[LoadQueue.scala 233:38:@9685.8]
  wire  _T_24863; // @[LoadQueue.scala 234:11:@9694.8]
  wire  _T_24864; // @[LoadQueue.scala 233:103:@9695.8]
  wire  _GEN_540; // @[LoadQueue.scala 230:110:@9676.6]
  wire  loadRequest_1; // @[LoadQueue.scala 229:71:@9670.4]
  wire [7:0] _T_24190; // @[Mux.scala 31:69:@9237.4]
  wire  _T_24780; // @[LoadQueue.scala 229:41:@9618.4]
  wire  _T_24781; // @[LoadQueue.scala 229:38:@9619.4]
  wire  _T_24783; // @[LoadQueue.scala 230:12:@9621.6]
  reg  prevPriorityRequest_0; // @[LoadQueue.scala 207:36:@9530.4]
  reg [31:0] _RAND_250;
  wire  _T_24785; // @[LoadQueue.scala 230:46:@9622.6]
  wire  _T_24786; // @[LoadQueue.scala 230:43:@9623.6]
  wire  _T_24788; // @[LoadQueue.scala 230:84:@9624.6]
  wire  _T_24789; // @[LoadQueue.scala 230:81:@9625.6]
  wire  _T_24792; // @[LoadQueue.scala 233:86:@9628.8]
  wire  _T_24793; // @[LoadQueue.scala 233:86:@9629.8]
  wire  _T_24794; // @[LoadQueue.scala 233:86:@9630.8]
  wire  _T_24795; // @[LoadQueue.scala 233:86:@9631.8]
  wire  _T_24796; // @[LoadQueue.scala 233:86:@9632.8]
  wire  _T_24797; // @[LoadQueue.scala 233:86:@9633.8]
  wire  _T_24798; // @[LoadQueue.scala 233:86:@9634.8]
  wire  _T_24800; // @[LoadQueue.scala 233:38:@9635.8]
  wire  _T_24811; // @[LoadQueue.scala 234:11:@9644.8]
  wire  _T_24812; // @[LoadQueue.scala 233:103:@9645.8]
  wire  _GEN_536; // @[LoadQueue.scala 230:110:@9626.6]
  wire  loadRequest_0; // @[LoadQueue.scala 229:71:@9620.4]
  wire [7:0] _T_24191; // @[Mux.scala 31:69:@9238.4]
  wire  _T_24192; // @[OneHot.scala 66:30:@9239.4]
  wire  _T_24193; // @[OneHot.scala 66:30:@9240.4]
  wire  _T_24194; // @[OneHot.scala 66:30:@9241.4]
  wire  _T_24195; // @[OneHot.scala 66:30:@9242.4]
  wire  _T_24196; // @[OneHot.scala 66:30:@9243.4]
  wire  _T_24197; // @[OneHot.scala 66:30:@9244.4]
  wire  _T_24198; // @[OneHot.scala 66:30:@9245.4]
  wire  _T_24199; // @[OneHot.scala 66:30:@9246.4]
  wire [7:0] _T_24224; // @[Mux.scala 31:69:@9256.4]
  wire [7:0] _T_24225; // @[Mux.scala 31:69:@9257.4]
  wire [7:0] _T_24226; // @[Mux.scala 31:69:@9258.4]
  wire [7:0] _T_24227; // @[Mux.scala 31:69:@9259.4]
  wire [7:0] _T_24228; // @[Mux.scala 31:69:@9260.4]
  wire [7:0] _T_24229; // @[Mux.scala 31:69:@9261.4]
  wire [7:0] _T_24230; // @[Mux.scala 31:69:@9262.4]
  wire [7:0] _T_24231; // @[Mux.scala 31:69:@9263.4]
  wire  _T_24232; // @[OneHot.scala 66:30:@9264.4]
  wire  _T_24233; // @[OneHot.scala 66:30:@9265.4]
  wire  _T_24234; // @[OneHot.scala 66:30:@9266.4]
  wire  _T_24235; // @[OneHot.scala 66:30:@9267.4]
  wire  _T_24236; // @[OneHot.scala 66:30:@9268.4]
  wire  _T_24237; // @[OneHot.scala 66:30:@9269.4]
  wire  _T_24238; // @[OneHot.scala 66:30:@9270.4]
  wire  _T_24239; // @[OneHot.scala 66:30:@9271.4]
  wire [7:0] _T_24264; // @[Mux.scala 31:69:@9281.4]
  wire [7:0] _T_24265; // @[Mux.scala 31:69:@9282.4]
  wire [7:0] _T_24266; // @[Mux.scala 31:69:@9283.4]
  wire [7:0] _T_24267; // @[Mux.scala 31:69:@9284.4]
  wire [7:0] _T_24268; // @[Mux.scala 31:69:@9285.4]
  wire [7:0] _T_24269; // @[Mux.scala 31:69:@9286.4]
  wire [7:0] _T_24270; // @[Mux.scala 31:69:@9287.4]
  wire [7:0] _T_24271; // @[Mux.scala 31:69:@9288.4]
  wire  _T_24272; // @[OneHot.scala 66:30:@9289.4]
  wire  _T_24273; // @[OneHot.scala 66:30:@9290.4]
  wire  _T_24274; // @[OneHot.scala 66:30:@9291.4]
  wire  _T_24275; // @[OneHot.scala 66:30:@9292.4]
  wire  _T_24276; // @[OneHot.scala 66:30:@9293.4]
  wire  _T_24277; // @[OneHot.scala 66:30:@9294.4]
  wire  _T_24278; // @[OneHot.scala 66:30:@9295.4]
  wire  _T_24279; // @[OneHot.scala 66:30:@9296.4]
  wire [7:0] _T_24304; // @[Mux.scala 31:69:@9306.4]
  wire [7:0] _T_24305; // @[Mux.scala 31:69:@9307.4]
  wire [7:0] _T_24306; // @[Mux.scala 31:69:@9308.4]
  wire [7:0] _T_24307; // @[Mux.scala 31:69:@9309.4]
  wire [7:0] _T_24308; // @[Mux.scala 31:69:@9310.4]
  wire [7:0] _T_24309; // @[Mux.scala 31:69:@9311.4]
  wire [7:0] _T_24310; // @[Mux.scala 31:69:@9312.4]
  wire [7:0] _T_24311; // @[Mux.scala 31:69:@9313.4]
  wire  _T_24312; // @[OneHot.scala 66:30:@9314.4]
  wire  _T_24313; // @[OneHot.scala 66:30:@9315.4]
  wire  _T_24314; // @[OneHot.scala 66:30:@9316.4]
  wire  _T_24315; // @[OneHot.scala 66:30:@9317.4]
  wire  _T_24316; // @[OneHot.scala 66:30:@9318.4]
  wire  _T_24317; // @[OneHot.scala 66:30:@9319.4]
  wire  _T_24318; // @[OneHot.scala 66:30:@9320.4]
  wire  _T_24319; // @[OneHot.scala 66:30:@9321.4]
  wire [7:0] _T_24344; // @[Mux.scala 31:69:@9331.4]
  wire [7:0] _T_24345; // @[Mux.scala 31:69:@9332.4]
  wire [7:0] _T_24346; // @[Mux.scala 31:69:@9333.4]
  wire [7:0] _T_24347; // @[Mux.scala 31:69:@9334.4]
  wire [7:0] _T_24348; // @[Mux.scala 31:69:@9335.4]
  wire [7:0] _T_24349; // @[Mux.scala 31:69:@9336.4]
  wire [7:0] _T_24350; // @[Mux.scala 31:69:@9337.4]
  wire [7:0] _T_24351; // @[Mux.scala 31:69:@9338.4]
  wire  _T_24352; // @[OneHot.scala 66:30:@9339.4]
  wire  _T_24353; // @[OneHot.scala 66:30:@9340.4]
  wire  _T_24354; // @[OneHot.scala 66:30:@9341.4]
  wire  _T_24355; // @[OneHot.scala 66:30:@9342.4]
  wire  _T_24356; // @[OneHot.scala 66:30:@9343.4]
  wire  _T_24357; // @[OneHot.scala 66:30:@9344.4]
  wire  _T_24358; // @[OneHot.scala 66:30:@9345.4]
  wire  _T_24359; // @[OneHot.scala 66:30:@9346.4]
  wire [7:0] _T_24384; // @[Mux.scala 31:69:@9356.4]
  wire [7:0] _T_24385; // @[Mux.scala 31:69:@9357.4]
  wire [7:0] _T_24386; // @[Mux.scala 31:69:@9358.4]
  wire [7:0] _T_24387; // @[Mux.scala 31:69:@9359.4]
  wire [7:0] _T_24388; // @[Mux.scala 31:69:@9360.4]
  wire [7:0] _T_24389; // @[Mux.scala 31:69:@9361.4]
  wire [7:0] _T_24390; // @[Mux.scala 31:69:@9362.4]
  wire [7:0] _T_24391; // @[Mux.scala 31:69:@9363.4]
  wire  _T_24392; // @[OneHot.scala 66:30:@9364.4]
  wire  _T_24393; // @[OneHot.scala 66:30:@9365.4]
  wire  _T_24394; // @[OneHot.scala 66:30:@9366.4]
  wire  _T_24395; // @[OneHot.scala 66:30:@9367.4]
  wire  _T_24396; // @[OneHot.scala 66:30:@9368.4]
  wire  _T_24397; // @[OneHot.scala 66:30:@9369.4]
  wire  _T_24398; // @[OneHot.scala 66:30:@9370.4]
  wire  _T_24399; // @[OneHot.scala 66:30:@9371.4]
  wire [7:0] _T_24424; // @[Mux.scala 31:69:@9381.4]
  wire [7:0] _T_24425; // @[Mux.scala 31:69:@9382.4]
  wire [7:0] _T_24426; // @[Mux.scala 31:69:@9383.4]
  wire [7:0] _T_24427; // @[Mux.scala 31:69:@9384.4]
  wire [7:0] _T_24428; // @[Mux.scala 31:69:@9385.4]
  wire [7:0] _T_24429; // @[Mux.scala 31:69:@9386.4]
  wire [7:0] _T_24430; // @[Mux.scala 31:69:@9387.4]
  wire [7:0] _T_24431; // @[Mux.scala 31:69:@9388.4]
  wire  _T_24432; // @[OneHot.scala 66:30:@9389.4]
  wire  _T_24433; // @[OneHot.scala 66:30:@9390.4]
  wire  _T_24434; // @[OneHot.scala 66:30:@9391.4]
  wire  _T_24435; // @[OneHot.scala 66:30:@9392.4]
  wire  _T_24436; // @[OneHot.scala 66:30:@9393.4]
  wire  _T_24437; // @[OneHot.scala 66:30:@9394.4]
  wire  _T_24438; // @[OneHot.scala 66:30:@9395.4]
  wire  _T_24439; // @[OneHot.scala 66:30:@9396.4]
  wire [7:0] _T_24464; // @[Mux.scala 31:69:@9406.4]
  wire [7:0] _T_24465; // @[Mux.scala 31:69:@9407.4]
  wire [7:0] _T_24466; // @[Mux.scala 31:69:@9408.4]
  wire [7:0] _T_24467; // @[Mux.scala 31:69:@9409.4]
  wire [7:0] _T_24468; // @[Mux.scala 31:69:@9410.4]
  wire [7:0] _T_24469; // @[Mux.scala 31:69:@9411.4]
  wire [7:0] _T_24470; // @[Mux.scala 31:69:@9412.4]
  wire [7:0] _T_24471; // @[Mux.scala 31:69:@9413.4]
  wire  _T_24472; // @[OneHot.scala 66:30:@9414.4]
  wire  _T_24473; // @[OneHot.scala 66:30:@9415.4]
  wire  _T_24474; // @[OneHot.scala 66:30:@9416.4]
  wire  _T_24475; // @[OneHot.scala 66:30:@9417.4]
  wire  _T_24476; // @[OneHot.scala 66:30:@9418.4]
  wire  _T_24477; // @[OneHot.scala 66:30:@9419.4]
  wire  _T_24478; // @[OneHot.scala 66:30:@9420.4]
  wire  _T_24479; // @[OneHot.scala 66:30:@9421.4]
  wire [7:0] _T_24520; // @[Mux.scala 19:72:@9437.4]
  wire [7:0] _T_24522; // @[Mux.scala 19:72:@9438.4]
  wire [7:0] _T_24529; // @[Mux.scala 19:72:@9445.4]
  wire [7:0] _T_24531; // @[Mux.scala 19:72:@9446.4]
  wire [7:0] _T_24538; // @[Mux.scala 19:72:@9453.4]
  wire [7:0] _T_24540; // @[Mux.scala 19:72:@9454.4]
  wire [7:0] _T_24547; // @[Mux.scala 19:72:@9461.4]
  wire [7:0] _T_24549; // @[Mux.scala 19:72:@9462.4]
  wire [7:0] _T_24556; // @[Mux.scala 19:72:@9469.4]
  wire [7:0] _T_24558; // @[Mux.scala 19:72:@9470.4]
  wire [7:0] _T_24565; // @[Mux.scala 19:72:@9477.4]
  wire [7:0] _T_24567; // @[Mux.scala 19:72:@9478.4]
  wire [7:0] _T_24574; // @[Mux.scala 19:72:@9485.4]
  wire [7:0] _T_24576; // @[Mux.scala 19:72:@9486.4]
  wire [7:0] _T_24583; // @[Mux.scala 19:72:@9493.4]
  wire [7:0] _T_24585; // @[Mux.scala 19:72:@9494.4]
  wire [7:0] _T_24586; // @[Mux.scala 19:72:@9495.4]
  wire [7:0] _T_24587; // @[Mux.scala 19:72:@9496.4]
  wire [7:0] _T_24588; // @[Mux.scala 19:72:@9497.4]
  wire [7:0] _T_24589; // @[Mux.scala 19:72:@9498.4]
  wire [7:0] _T_24590; // @[Mux.scala 19:72:@9499.4]
  wire [7:0] _T_24591; // @[Mux.scala 19:72:@9500.4]
  wire [7:0] _T_24592; // @[Mux.scala 19:72:@9501.4]
  wire  priorityLoadRequest_0; // @[Mux.scala 19:72:@9505.4]
  wire  priorityLoadRequest_1; // @[Mux.scala 19:72:@9507.4]
  wire  priorityLoadRequest_2; // @[Mux.scala 19:72:@9509.4]
  wire  priorityLoadRequest_3; // @[Mux.scala 19:72:@9511.4]
  wire  priorityLoadRequest_4; // @[Mux.scala 19:72:@9513.4]
  wire  priorityLoadRequest_5; // @[Mux.scala 19:72:@9515.4]
  wire  priorityLoadRequest_6; // @[Mux.scala 19:72:@9517.4]
  wire  priorityLoadRequest_7; // @[Mux.scala 19:72:@9519.4]
  wire  _GEN_512; // @[LoadQueue.scala 208:31:@9531.4]
  wire  _GEN_513; // @[LoadQueue.scala 208:31:@9531.4]
  wire  _GEN_514; // @[LoadQueue.scala 208:31:@9531.4]
  wire  _GEN_515; // @[LoadQueue.scala 208:31:@9531.4]
  wire  _GEN_516; // @[LoadQueue.scala 208:31:@9531.4]
  wire  _GEN_517; // @[LoadQueue.scala 208:31:@9531.4]
  wire  _GEN_518; // @[LoadQueue.scala 208:31:@9531.4]
  wire  _GEN_519; // @[LoadQueue.scala 208:31:@9531.4]
  wire [7:0] _T_24819; // @[LoadQueue.scala 238:58:@9653.8]
  wire [7:0] _T_24826; // @[LoadQueue.scala 238:96:@9660.8]
  wire  _T_24827; // @[LoadQueue.scala 238:61:@9661.8]
  wire  _T_24828; // @[LoadQueue.scala 237:64:@9662.8]
  wire  _GEN_537; // @[LoadQueue.scala 230:110:@9626.6]
  wire  bypassRequest_0; // @[LoadQueue.scala 229:71:@9620.4]
  wire  _GEN_520; // @[LoadQueue.scala 217:34:@9564.6]
  wire  _GEN_521; // @[LoadQueue.scala 215:23:@9560.4]
  wire [7:0] _T_24871; // @[LoadQueue.scala 238:58:@9703.8]
  wire [7:0] _T_24878; // @[LoadQueue.scala 238:96:@9710.8]
  wire  _T_24879; // @[LoadQueue.scala 238:61:@9711.8]
  wire  _T_24880; // @[LoadQueue.scala 237:64:@9712.8]
  wire  _GEN_541; // @[LoadQueue.scala 230:110:@9676.6]
  wire  bypassRequest_1; // @[LoadQueue.scala 229:71:@9670.4]
  wire  _GEN_522; // @[LoadQueue.scala 217:34:@9571.6]
  wire  _GEN_523; // @[LoadQueue.scala 215:23:@9567.4]
  wire [7:0] _T_24923; // @[LoadQueue.scala 238:58:@9753.8]
  wire [7:0] _T_24930; // @[LoadQueue.scala 238:96:@9760.8]
  wire  _T_24931; // @[LoadQueue.scala 238:61:@9761.8]
  wire  _T_24932; // @[LoadQueue.scala 237:64:@9762.8]
  wire  _GEN_545; // @[LoadQueue.scala 230:110:@9726.6]
  wire  bypassRequest_2; // @[LoadQueue.scala 229:71:@9720.4]
  wire  _GEN_524; // @[LoadQueue.scala 217:34:@9578.6]
  wire  _GEN_525; // @[LoadQueue.scala 215:23:@9574.4]
  wire [7:0] _T_24975; // @[LoadQueue.scala 238:58:@9803.8]
  wire [7:0] _T_24982; // @[LoadQueue.scala 238:96:@9810.8]
  wire  _T_24983; // @[LoadQueue.scala 238:61:@9811.8]
  wire  _T_24984; // @[LoadQueue.scala 237:64:@9812.8]
  wire  _GEN_549; // @[LoadQueue.scala 230:110:@9776.6]
  wire  bypassRequest_3; // @[LoadQueue.scala 229:71:@9770.4]
  wire  _GEN_526; // @[LoadQueue.scala 217:34:@9585.6]
  wire  _GEN_527; // @[LoadQueue.scala 215:23:@9581.4]
  wire [7:0] _T_25027; // @[LoadQueue.scala 238:58:@9853.8]
  wire [7:0] _T_25034; // @[LoadQueue.scala 238:96:@9860.8]
  wire  _T_25035; // @[LoadQueue.scala 238:61:@9861.8]
  wire  _T_25036; // @[LoadQueue.scala 237:64:@9862.8]
  wire  _GEN_553; // @[LoadQueue.scala 230:110:@9826.6]
  wire  bypassRequest_4; // @[LoadQueue.scala 229:71:@9820.4]
  wire  _GEN_528; // @[LoadQueue.scala 217:34:@9592.6]
  wire  _GEN_529; // @[LoadQueue.scala 215:23:@9588.4]
  wire [7:0] _T_25079; // @[LoadQueue.scala 238:58:@9903.8]
  wire [7:0] _T_25086; // @[LoadQueue.scala 238:96:@9910.8]
  wire  _T_25087; // @[LoadQueue.scala 238:61:@9911.8]
  wire  _T_25088; // @[LoadQueue.scala 237:64:@9912.8]
  wire  _GEN_557; // @[LoadQueue.scala 230:110:@9876.6]
  wire  bypassRequest_5; // @[LoadQueue.scala 229:71:@9870.4]
  wire  _GEN_530; // @[LoadQueue.scala 217:34:@9599.6]
  wire  _GEN_531; // @[LoadQueue.scala 215:23:@9595.4]
  wire [7:0] _T_25131; // @[LoadQueue.scala 238:58:@9953.8]
  wire [7:0] _T_25138; // @[LoadQueue.scala 238:96:@9960.8]
  wire  _T_25139; // @[LoadQueue.scala 238:61:@9961.8]
  wire  _T_25140; // @[LoadQueue.scala 237:64:@9962.8]
  wire  _GEN_561; // @[LoadQueue.scala 230:110:@9926.6]
  wire  bypassRequest_6; // @[LoadQueue.scala 229:71:@9920.4]
  wire  _GEN_532; // @[LoadQueue.scala 217:34:@9606.6]
  wire  _GEN_533; // @[LoadQueue.scala 215:23:@9602.4]
  wire [7:0] _T_25183; // @[LoadQueue.scala 238:58:@10003.8]
  wire [7:0] _T_25190; // @[LoadQueue.scala 238:96:@10010.8]
  wire  _T_25191; // @[LoadQueue.scala 238:61:@10011.8]
  wire  _T_25192; // @[LoadQueue.scala 237:64:@10012.8]
  wire  _GEN_565; // @[LoadQueue.scala 230:110:@9976.6]
  wire  bypassRequest_7; // @[LoadQueue.scala 229:71:@9970.4]
  wire  _GEN_534; // @[LoadQueue.scala 217:34:@9613.6]
  wire  _GEN_535; // @[LoadQueue.scala 215:23:@9609.4]
  wire  _T_25196; // @[LoadQueue.scala 247:28:@10018.4]
  wire  _T_25197; // @[LoadQueue.scala 247:28:@10019.4]
  wire  _T_25198; // @[LoadQueue.scala 247:28:@10020.4]
  wire  _T_25199; // @[LoadQueue.scala 247:28:@10021.4]
  wire  _T_25200; // @[LoadQueue.scala 247:28:@10022.4]
  wire  _T_25201; // @[LoadQueue.scala 247:28:@10023.4]
  wire  _T_25202; // @[LoadQueue.scala 247:28:@10024.4]
  wire [2:0] _T_25211; // @[Mux.scala 31:69:@10026.6]
  wire [2:0] _T_25212; // @[Mux.scala 31:69:@10027.6]
  wire [2:0] _T_25213; // @[Mux.scala 31:69:@10028.6]
  wire [2:0] _T_25214; // @[Mux.scala 31:69:@10029.6]
  wire [2:0] _T_25215; // @[Mux.scala 31:69:@10030.6]
  wire [2:0] _T_25216; // @[Mux.scala 31:69:@10031.6]
  wire [2:0] _T_25217; // @[Mux.scala 31:69:@10032.6]
  wire [31:0] _GEN_569; // @[LoadQueue.scala 248:24:@10033.6]
  wire [31:0] _GEN_570; // @[LoadQueue.scala 248:24:@10033.6]
  wire [31:0] _GEN_571; // @[LoadQueue.scala 248:24:@10033.6]
  wire [31:0] _GEN_572; // @[LoadQueue.scala 248:24:@10033.6]
  wire [31:0] _GEN_573; // @[LoadQueue.scala 248:24:@10033.6]
  wire [31:0] _GEN_574; // @[LoadQueue.scala 248:24:@10033.6]
  wire [31:0] _GEN_575; // @[LoadQueue.scala 248:24:@10033.6]
  wire  _T_25225; // @[LoadQueue.scala 261:41:@10044.6]
  wire  _GEN_578; // @[LoadQueue.scala 261:62:@10045.6]
  wire  _GEN_579; // @[LoadQueue.scala 259:25:@10040.4]
  wire  _T_25228; // @[LoadQueue.scala 261:41:@10052.6]
  wire  _GEN_580; // @[LoadQueue.scala 261:62:@10053.6]
  wire  _GEN_581; // @[LoadQueue.scala 259:25:@10048.4]
  wire  _T_25231; // @[LoadQueue.scala 261:41:@10060.6]
  wire  _GEN_582; // @[LoadQueue.scala 261:62:@10061.6]
  wire  _GEN_583; // @[LoadQueue.scala 259:25:@10056.4]
  wire  _T_25234; // @[LoadQueue.scala 261:41:@10068.6]
  wire  _GEN_584; // @[LoadQueue.scala 261:62:@10069.6]
  wire  _GEN_585; // @[LoadQueue.scala 259:25:@10064.4]
  wire  _T_25237; // @[LoadQueue.scala 261:41:@10076.6]
  wire  _GEN_586; // @[LoadQueue.scala 261:62:@10077.6]
  wire  _GEN_587; // @[LoadQueue.scala 259:25:@10072.4]
  wire  _T_25240; // @[LoadQueue.scala 261:41:@10084.6]
  wire  _GEN_588; // @[LoadQueue.scala 261:62:@10085.6]
  wire  _GEN_589; // @[LoadQueue.scala 259:25:@10080.4]
  wire  _T_25243; // @[LoadQueue.scala 261:41:@10092.6]
  wire  _GEN_590; // @[LoadQueue.scala 261:62:@10093.6]
  wire  _GEN_591; // @[LoadQueue.scala 259:25:@10088.4]
  wire  _T_25246; // @[LoadQueue.scala 261:41:@10100.6]
  wire  _GEN_592; // @[LoadQueue.scala 261:62:@10101.6]
  wire  _GEN_593; // @[LoadQueue.scala 259:25:@10096.4]
  wire [31:0] _GEN_594; // @[LoadQueue.scala 269:44:@10108.6]
  wire [31:0] _GEN_595; // @[LoadQueue.scala 267:32:@10104.4]
  wire [31:0] _GEN_596; // @[LoadQueue.scala 269:44:@10115.6]
  wire [31:0] _GEN_597; // @[LoadQueue.scala 267:32:@10111.4]
  wire [31:0] _GEN_598; // @[LoadQueue.scala 269:44:@10122.6]
  wire [31:0] _GEN_599; // @[LoadQueue.scala 267:32:@10118.4]
  wire [31:0] _GEN_600; // @[LoadQueue.scala 269:44:@10129.6]
  wire [31:0] _GEN_601; // @[LoadQueue.scala 267:32:@10125.4]
  wire [31:0] _GEN_602; // @[LoadQueue.scala 269:44:@10136.6]
  wire [31:0] _GEN_603; // @[LoadQueue.scala 267:32:@10132.4]
  wire [31:0] _GEN_604; // @[LoadQueue.scala 269:44:@10143.6]
  wire [31:0] _GEN_605; // @[LoadQueue.scala 267:32:@10139.4]
  wire [31:0] _GEN_606; // @[LoadQueue.scala 269:44:@10150.6]
  wire [31:0] _GEN_607; // @[LoadQueue.scala 267:32:@10146.4]
  wire [31:0] _GEN_608; // @[LoadQueue.scala 269:44:@10157.6]
  wire [31:0] _GEN_609; // @[LoadQueue.scala 267:32:@10153.4]
  wire  entriesPorts_0_0; // @[LoadQueue.scala 286:69:@10161.4]
  wire  entriesPorts_0_1; // @[LoadQueue.scala 286:69:@10163.4]
  wire  entriesPorts_0_2; // @[LoadQueue.scala 286:69:@10165.4]
  wire  entriesPorts_0_3; // @[LoadQueue.scala 286:69:@10167.4]
  wire  entriesPorts_0_4; // @[LoadQueue.scala 286:69:@10169.4]
  wire  entriesPorts_0_5; // @[LoadQueue.scala 286:69:@10171.4]
  wire  entriesPorts_0_6; // @[LoadQueue.scala 286:69:@10173.4]
  wire  entriesPorts_0_7; // @[LoadQueue.scala 286:69:@10175.4]
  wire  _T_25659; // @[LoadQueue.scala 298:86:@10195.4]
  wire  _T_25660; // @[LoadQueue.scala 298:83:@10196.4]
  wire  _T_25662; // @[LoadQueue.scala 298:86:@10197.4]
  wire  _T_25663; // @[LoadQueue.scala 298:83:@10198.4]
  wire  _T_25665; // @[LoadQueue.scala 298:86:@10199.4]
  wire  _T_25666; // @[LoadQueue.scala 298:83:@10200.4]
  wire  _T_25668; // @[LoadQueue.scala 298:86:@10201.4]
  wire  _T_25669; // @[LoadQueue.scala 298:83:@10202.4]
  wire  _T_25671; // @[LoadQueue.scala 298:86:@10203.4]
  wire  _T_25672; // @[LoadQueue.scala 298:83:@10204.4]
  wire  _T_25674; // @[LoadQueue.scala 298:86:@10205.4]
  wire  _T_25675; // @[LoadQueue.scala 298:83:@10206.4]
  wire  _T_25677; // @[LoadQueue.scala 298:86:@10207.4]
  wire  _T_25678; // @[LoadQueue.scala 298:83:@10208.4]
  wire  _T_25680; // @[LoadQueue.scala 298:86:@10209.4]
  wire  _T_25681; // @[LoadQueue.scala 298:83:@10210.4]
  wire [7:0] _T_25732; // @[Mux.scala 31:69:@10240.4]
  wire [7:0] _T_25733; // @[Mux.scala 31:69:@10241.4]
  wire [7:0] _T_25734; // @[Mux.scala 31:69:@10242.4]
  wire [7:0] _T_25735; // @[Mux.scala 31:69:@10243.4]
  wire [7:0] _T_25736; // @[Mux.scala 31:69:@10244.4]
  wire [7:0] _T_25737; // @[Mux.scala 31:69:@10245.4]
  wire [7:0] _T_25738; // @[Mux.scala 31:69:@10246.4]
  wire [7:0] _T_25739; // @[Mux.scala 31:69:@10247.4]
  wire  _T_25740; // @[OneHot.scala 66:30:@10248.4]
  wire  _T_25741; // @[OneHot.scala 66:30:@10249.4]
  wire  _T_25742; // @[OneHot.scala 66:30:@10250.4]
  wire  _T_25743; // @[OneHot.scala 66:30:@10251.4]
  wire  _T_25744; // @[OneHot.scala 66:30:@10252.4]
  wire  _T_25745; // @[OneHot.scala 66:30:@10253.4]
  wire  _T_25746; // @[OneHot.scala 66:30:@10254.4]
  wire  _T_25747; // @[OneHot.scala 66:30:@10255.4]
  wire [7:0] _T_25772; // @[Mux.scala 31:69:@10265.4]
  wire [7:0] _T_25773; // @[Mux.scala 31:69:@10266.4]
  wire [7:0] _T_25774; // @[Mux.scala 31:69:@10267.4]
  wire [7:0] _T_25775; // @[Mux.scala 31:69:@10268.4]
  wire [7:0] _T_25776; // @[Mux.scala 31:69:@10269.4]
  wire [7:0] _T_25777; // @[Mux.scala 31:69:@10270.4]
  wire [7:0] _T_25778; // @[Mux.scala 31:69:@10271.4]
  wire [7:0] _T_25779; // @[Mux.scala 31:69:@10272.4]
  wire  _T_25780; // @[OneHot.scala 66:30:@10273.4]
  wire  _T_25781; // @[OneHot.scala 66:30:@10274.4]
  wire  _T_25782; // @[OneHot.scala 66:30:@10275.4]
  wire  _T_25783; // @[OneHot.scala 66:30:@10276.4]
  wire  _T_25784; // @[OneHot.scala 66:30:@10277.4]
  wire  _T_25785; // @[OneHot.scala 66:30:@10278.4]
  wire  _T_25786; // @[OneHot.scala 66:30:@10279.4]
  wire  _T_25787; // @[OneHot.scala 66:30:@10280.4]
  wire [7:0] _T_25812; // @[Mux.scala 31:69:@10290.4]
  wire [7:0] _T_25813; // @[Mux.scala 31:69:@10291.4]
  wire [7:0] _T_25814; // @[Mux.scala 31:69:@10292.4]
  wire [7:0] _T_25815; // @[Mux.scala 31:69:@10293.4]
  wire [7:0] _T_25816; // @[Mux.scala 31:69:@10294.4]
  wire [7:0] _T_25817; // @[Mux.scala 31:69:@10295.4]
  wire [7:0] _T_25818; // @[Mux.scala 31:69:@10296.4]
  wire [7:0] _T_25819; // @[Mux.scala 31:69:@10297.4]
  wire  _T_25820; // @[OneHot.scala 66:30:@10298.4]
  wire  _T_25821; // @[OneHot.scala 66:30:@10299.4]
  wire  _T_25822; // @[OneHot.scala 66:30:@10300.4]
  wire  _T_25823; // @[OneHot.scala 66:30:@10301.4]
  wire  _T_25824; // @[OneHot.scala 66:30:@10302.4]
  wire  _T_25825; // @[OneHot.scala 66:30:@10303.4]
  wire  _T_25826; // @[OneHot.scala 66:30:@10304.4]
  wire  _T_25827; // @[OneHot.scala 66:30:@10305.4]
  wire [7:0] _T_25852; // @[Mux.scala 31:69:@10315.4]
  wire [7:0] _T_25853; // @[Mux.scala 31:69:@10316.4]
  wire [7:0] _T_25854; // @[Mux.scala 31:69:@10317.4]
  wire [7:0] _T_25855; // @[Mux.scala 31:69:@10318.4]
  wire [7:0] _T_25856; // @[Mux.scala 31:69:@10319.4]
  wire [7:0] _T_25857; // @[Mux.scala 31:69:@10320.4]
  wire [7:0] _T_25858; // @[Mux.scala 31:69:@10321.4]
  wire [7:0] _T_25859; // @[Mux.scala 31:69:@10322.4]
  wire  _T_25860; // @[OneHot.scala 66:30:@10323.4]
  wire  _T_25861; // @[OneHot.scala 66:30:@10324.4]
  wire  _T_25862; // @[OneHot.scala 66:30:@10325.4]
  wire  _T_25863; // @[OneHot.scala 66:30:@10326.4]
  wire  _T_25864; // @[OneHot.scala 66:30:@10327.4]
  wire  _T_25865; // @[OneHot.scala 66:30:@10328.4]
  wire  _T_25866; // @[OneHot.scala 66:30:@10329.4]
  wire  _T_25867; // @[OneHot.scala 66:30:@10330.4]
  wire [7:0] _T_25892; // @[Mux.scala 31:69:@10340.4]
  wire [7:0] _T_25893; // @[Mux.scala 31:69:@10341.4]
  wire [7:0] _T_25894; // @[Mux.scala 31:69:@10342.4]
  wire [7:0] _T_25895; // @[Mux.scala 31:69:@10343.4]
  wire [7:0] _T_25896; // @[Mux.scala 31:69:@10344.4]
  wire [7:0] _T_25897; // @[Mux.scala 31:69:@10345.4]
  wire [7:0] _T_25898; // @[Mux.scala 31:69:@10346.4]
  wire [7:0] _T_25899; // @[Mux.scala 31:69:@10347.4]
  wire  _T_25900; // @[OneHot.scala 66:30:@10348.4]
  wire  _T_25901; // @[OneHot.scala 66:30:@10349.4]
  wire  _T_25902; // @[OneHot.scala 66:30:@10350.4]
  wire  _T_25903; // @[OneHot.scala 66:30:@10351.4]
  wire  _T_25904; // @[OneHot.scala 66:30:@10352.4]
  wire  _T_25905; // @[OneHot.scala 66:30:@10353.4]
  wire  _T_25906; // @[OneHot.scala 66:30:@10354.4]
  wire  _T_25907; // @[OneHot.scala 66:30:@10355.4]
  wire [7:0] _T_25932; // @[Mux.scala 31:69:@10365.4]
  wire [7:0] _T_25933; // @[Mux.scala 31:69:@10366.4]
  wire [7:0] _T_25934; // @[Mux.scala 31:69:@10367.4]
  wire [7:0] _T_25935; // @[Mux.scala 31:69:@10368.4]
  wire [7:0] _T_25936; // @[Mux.scala 31:69:@10369.4]
  wire [7:0] _T_25937; // @[Mux.scala 31:69:@10370.4]
  wire [7:0] _T_25938; // @[Mux.scala 31:69:@10371.4]
  wire [7:0] _T_25939; // @[Mux.scala 31:69:@10372.4]
  wire  _T_25940; // @[OneHot.scala 66:30:@10373.4]
  wire  _T_25941; // @[OneHot.scala 66:30:@10374.4]
  wire  _T_25942; // @[OneHot.scala 66:30:@10375.4]
  wire  _T_25943; // @[OneHot.scala 66:30:@10376.4]
  wire  _T_25944; // @[OneHot.scala 66:30:@10377.4]
  wire  _T_25945; // @[OneHot.scala 66:30:@10378.4]
  wire  _T_25946; // @[OneHot.scala 66:30:@10379.4]
  wire  _T_25947; // @[OneHot.scala 66:30:@10380.4]
  wire [7:0] _T_25972; // @[Mux.scala 31:69:@10390.4]
  wire [7:0] _T_25973; // @[Mux.scala 31:69:@10391.4]
  wire [7:0] _T_25974; // @[Mux.scala 31:69:@10392.4]
  wire [7:0] _T_25975; // @[Mux.scala 31:69:@10393.4]
  wire [7:0] _T_25976; // @[Mux.scala 31:69:@10394.4]
  wire [7:0] _T_25977; // @[Mux.scala 31:69:@10395.4]
  wire [7:0] _T_25978; // @[Mux.scala 31:69:@10396.4]
  wire [7:0] _T_25979; // @[Mux.scala 31:69:@10397.4]
  wire  _T_25980; // @[OneHot.scala 66:30:@10398.4]
  wire  _T_25981; // @[OneHot.scala 66:30:@10399.4]
  wire  _T_25982; // @[OneHot.scala 66:30:@10400.4]
  wire  _T_25983; // @[OneHot.scala 66:30:@10401.4]
  wire  _T_25984; // @[OneHot.scala 66:30:@10402.4]
  wire  _T_25985; // @[OneHot.scala 66:30:@10403.4]
  wire  _T_25986; // @[OneHot.scala 66:30:@10404.4]
  wire  _T_25987; // @[OneHot.scala 66:30:@10405.4]
  wire [7:0] _T_26012; // @[Mux.scala 31:69:@10415.4]
  wire [7:0] _T_26013; // @[Mux.scala 31:69:@10416.4]
  wire [7:0] _T_26014; // @[Mux.scala 31:69:@10417.4]
  wire [7:0] _T_26015; // @[Mux.scala 31:69:@10418.4]
  wire [7:0] _T_26016; // @[Mux.scala 31:69:@10419.4]
  wire [7:0] _T_26017; // @[Mux.scala 31:69:@10420.4]
  wire [7:0] _T_26018; // @[Mux.scala 31:69:@10421.4]
  wire [7:0] _T_26019; // @[Mux.scala 31:69:@10422.4]
  wire  _T_26020; // @[OneHot.scala 66:30:@10423.4]
  wire  _T_26021; // @[OneHot.scala 66:30:@10424.4]
  wire  _T_26022; // @[OneHot.scala 66:30:@10425.4]
  wire  _T_26023; // @[OneHot.scala 66:30:@10426.4]
  wire  _T_26024; // @[OneHot.scala 66:30:@10427.4]
  wire  _T_26025; // @[OneHot.scala 66:30:@10428.4]
  wire  _T_26026; // @[OneHot.scala 66:30:@10429.4]
  wire  _T_26027; // @[OneHot.scala 66:30:@10430.4]
  wire [7:0] _T_26068; // @[Mux.scala 19:72:@10446.4]
  wire [7:0] _T_26070; // @[Mux.scala 19:72:@10447.4]
  wire [7:0] _T_26077; // @[Mux.scala 19:72:@10454.4]
  wire [7:0] _T_26079; // @[Mux.scala 19:72:@10455.4]
  wire [7:0] _T_26086; // @[Mux.scala 19:72:@10462.4]
  wire [7:0] _T_26088; // @[Mux.scala 19:72:@10463.4]
  wire [7:0] _T_26095; // @[Mux.scala 19:72:@10470.4]
  wire [7:0] _T_26097; // @[Mux.scala 19:72:@10471.4]
  wire [7:0] _T_26104; // @[Mux.scala 19:72:@10478.4]
  wire [7:0] _T_26106; // @[Mux.scala 19:72:@10479.4]
  wire [7:0] _T_26113; // @[Mux.scala 19:72:@10486.4]
  wire [7:0] _T_26115; // @[Mux.scala 19:72:@10487.4]
  wire [7:0] _T_26122; // @[Mux.scala 19:72:@10494.4]
  wire [7:0] _T_26124; // @[Mux.scala 19:72:@10495.4]
  wire [7:0] _T_26131; // @[Mux.scala 19:72:@10502.4]
  wire [7:0] _T_26133; // @[Mux.scala 19:72:@10503.4]
  wire [7:0] _T_26134; // @[Mux.scala 19:72:@10504.4]
  wire [7:0] _T_26135; // @[Mux.scala 19:72:@10505.4]
  wire [7:0] _T_26136; // @[Mux.scala 19:72:@10506.4]
  wire [7:0] _T_26137; // @[Mux.scala 19:72:@10507.4]
  wire [7:0] _T_26138; // @[Mux.scala 19:72:@10508.4]
  wire [7:0] _T_26139; // @[Mux.scala 19:72:@10509.4]
  wire [7:0] _T_26140; // @[Mux.scala 19:72:@10510.4]
  wire  inputPriorityPorts_0_0; // @[Mux.scala 19:72:@10514.4]
  wire  inputPriorityPorts_0_1; // @[Mux.scala 19:72:@10516.4]
  wire  inputPriorityPorts_0_2; // @[Mux.scala 19:72:@10518.4]
  wire  inputPriorityPorts_0_3; // @[Mux.scala 19:72:@10520.4]
  wire  inputPriorityPorts_0_4; // @[Mux.scala 19:72:@10522.4]
  wire  inputPriorityPorts_0_5; // @[Mux.scala 19:72:@10524.4]
  wire  inputPriorityPorts_0_6; // @[Mux.scala 19:72:@10526.4]
  wire  inputPriorityPorts_0_7; // @[Mux.scala 19:72:@10528.4]
  wire [7:0] _T_26254; // @[Mux.scala 31:69:@10558.4]
  wire [7:0] _T_26255; // @[Mux.scala 31:69:@10559.4]
  wire [7:0] _T_26256; // @[Mux.scala 31:69:@10560.4]
  wire [7:0] _T_26257; // @[Mux.scala 31:69:@10561.4]
  wire [7:0] _T_26258; // @[Mux.scala 31:69:@10562.4]
  wire [7:0] _T_26259; // @[Mux.scala 31:69:@10563.4]
  wire [7:0] _T_26260; // @[Mux.scala 31:69:@10564.4]
  wire [7:0] _T_26261; // @[Mux.scala 31:69:@10565.4]
  wire  _T_26262; // @[OneHot.scala 66:30:@10566.4]
  wire  _T_26263; // @[OneHot.scala 66:30:@10567.4]
  wire  _T_26264; // @[OneHot.scala 66:30:@10568.4]
  wire  _T_26265; // @[OneHot.scala 66:30:@10569.4]
  wire  _T_26266; // @[OneHot.scala 66:30:@10570.4]
  wire  _T_26267; // @[OneHot.scala 66:30:@10571.4]
  wire  _T_26268; // @[OneHot.scala 66:30:@10572.4]
  wire  _T_26269; // @[OneHot.scala 66:30:@10573.4]
  wire [7:0] _T_26294; // @[Mux.scala 31:69:@10583.4]
  wire [7:0] _T_26295; // @[Mux.scala 31:69:@10584.4]
  wire [7:0] _T_26296; // @[Mux.scala 31:69:@10585.4]
  wire [7:0] _T_26297; // @[Mux.scala 31:69:@10586.4]
  wire [7:0] _T_26298; // @[Mux.scala 31:69:@10587.4]
  wire [7:0] _T_26299; // @[Mux.scala 31:69:@10588.4]
  wire [7:0] _T_26300; // @[Mux.scala 31:69:@10589.4]
  wire [7:0] _T_26301; // @[Mux.scala 31:69:@10590.4]
  wire  _T_26302; // @[OneHot.scala 66:30:@10591.4]
  wire  _T_26303; // @[OneHot.scala 66:30:@10592.4]
  wire  _T_26304; // @[OneHot.scala 66:30:@10593.4]
  wire  _T_26305; // @[OneHot.scala 66:30:@10594.4]
  wire  _T_26306; // @[OneHot.scala 66:30:@10595.4]
  wire  _T_26307; // @[OneHot.scala 66:30:@10596.4]
  wire  _T_26308; // @[OneHot.scala 66:30:@10597.4]
  wire  _T_26309; // @[OneHot.scala 66:30:@10598.4]
  wire [7:0] _T_26334; // @[Mux.scala 31:69:@10608.4]
  wire [7:0] _T_26335; // @[Mux.scala 31:69:@10609.4]
  wire [7:0] _T_26336; // @[Mux.scala 31:69:@10610.4]
  wire [7:0] _T_26337; // @[Mux.scala 31:69:@10611.4]
  wire [7:0] _T_26338; // @[Mux.scala 31:69:@10612.4]
  wire [7:0] _T_26339; // @[Mux.scala 31:69:@10613.4]
  wire [7:0] _T_26340; // @[Mux.scala 31:69:@10614.4]
  wire [7:0] _T_26341; // @[Mux.scala 31:69:@10615.4]
  wire  _T_26342; // @[OneHot.scala 66:30:@10616.4]
  wire  _T_26343; // @[OneHot.scala 66:30:@10617.4]
  wire  _T_26344; // @[OneHot.scala 66:30:@10618.4]
  wire  _T_26345; // @[OneHot.scala 66:30:@10619.4]
  wire  _T_26346; // @[OneHot.scala 66:30:@10620.4]
  wire  _T_26347; // @[OneHot.scala 66:30:@10621.4]
  wire  _T_26348; // @[OneHot.scala 66:30:@10622.4]
  wire  _T_26349; // @[OneHot.scala 66:30:@10623.4]
  wire [7:0] _T_26374; // @[Mux.scala 31:69:@10633.4]
  wire [7:0] _T_26375; // @[Mux.scala 31:69:@10634.4]
  wire [7:0] _T_26376; // @[Mux.scala 31:69:@10635.4]
  wire [7:0] _T_26377; // @[Mux.scala 31:69:@10636.4]
  wire [7:0] _T_26378; // @[Mux.scala 31:69:@10637.4]
  wire [7:0] _T_26379; // @[Mux.scala 31:69:@10638.4]
  wire [7:0] _T_26380; // @[Mux.scala 31:69:@10639.4]
  wire [7:0] _T_26381; // @[Mux.scala 31:69:@10640.4]
  wire  _T_26382; // @[OneHot.scala 66:30:@10641.4]
  wire  _T_26383; // @[OneHot.scala 66:30:@10642.4]
  wire  _T_26384; // @[OneHot.scala 66:30:@10643.4]
  wire  _T_26385; // @[OneHot.scala 66:30:@10644.4]
  wire  _T_26386; // @[OneHot.scala 66:30:@10645.4]
  wire  _T_26387; // @[OneHot.scala 66:30:@10646.4]
  wire  _T_26388; // @[OneHot.scala 66:30:@10647.4]
  wire  _T_26389; // @[OneHot.scala 66:30:@10648.4]
  wire [7:0] _T_26414; // @[Mux.scala 31:69:@10658.4]
  wire [7:0] _T_26415; // @[Mux.scala 31:69:@10659.4]
  wire [7:0] _T_26416; // @[Mux.scala 31:69:@10660.4]
  wire [7:0] _T_26417; // @[Mux.scala 31:69:@10661.4]
  wire [7:0] _T_26418; // @[Mux.scala 31:69:@10662.4]
  wire [7:0] _T_26419; // @[Mux.scala 31:69:@10663.4]
  wire [7:0] _T_26420; // @[Mux.scala 31:69:@10664.4]
  wire [7:0] _T_26421; // @[Mux.scala 31:69:@10665.4]
  wire  _T_26422; // @[OneHot.scala 66:30:@10666.4]
  wire  _T_26423; // @[OneHot.scala 66:30:@10667.4]
  wire  _T_26424; // @[OneHot.scala 66:30:@10668.4]
  wire  _T_26425; // @[OneHot.scala 66:30:@10669.4]
  wire  _T_26426; // @[OneHot.scala 66:30:@10670.4]
  wire  _T_26427; // @[OneHot.scala 66:30:@10671.4]
  wire  _T_26428; // @[OneHot.scala 66:30:@10672.4]
  wire  _T_26429; // @[OneHot.scala 66:30:@10673.4]
  wire [7:0] _T_26454; // @[Mux.scala 31:69:@10683.4]
  wire [7:0] _T_26455; // @[Mux.scala 31:69:@10684.4]
  wire [7:0] _T_26456; // @[Mux.scala 31:69:@10685.4]
  wire [7:0] _T_26457; // @[Mux.scala 31:69:@10686.4]
  wire [7:0] _T_26458; // @[Mux.scala 31:69:@10687.4]
  wire [7:0] _T_26459; // @[Mux.scala 31:69:@10688.4]
  wire [7:0] _T_26460; // @[Mux.scala 31:69:@10689.4]
  wire [7:0] _T_26461; // @[Mux.scala 31:69:@10690.4]
  wire  _T_26462; // @[OneHot.scala 66:30:@10691.4]
  wire  _T_26463; // @[OneHot.scala 66:30:@10692.4]
  wire  _T_26464; // @[OneHot.scala 66:30:@10693.4]
  wire  _T_26465; // @[OneHot.scala 66:30:@10694.4]
  wire  _T_26466; // @[OneHot.scala 66:30:@10695.4]
  wire  _T_26467; // @[OneHot.scala 66:30:@10696.4]
  wire  _T_26468; // @[OneHot.scala 66:30:@10697.4]
  wire  _T_26469; // @[OneHot.scala 66:30:@10698.4]
  wire [7:0] _T_26494; // @[Mux.scala 31:69:@10708.4]
  wire [7:0] _T_26495; // @[Mux.scala 31:69:@10709.4]
  wire [7:0] _T_26496; // @[Mux.scala 31:69:@10710.4]
  wire [7:0] _T_26497; // @[Mux.scala 31:69:@10711.4]
  wire [7:0] _T_26498; // @[Mux.scala 31:69:@10712.4]
  wire [7:0] _T_26499; // @[Mux.scala 31:69:@10713.4]
  wire [7:0] _T_26500; // @[Mux.scala 31:69:@10714.4]
  wire [7:0] _T_26501; // @[Mux.scala 31:69:@10715.4]
  wire  _T_26502; // @[OneHot.scala 66:30:@10716.4]
  wire  _T_26503; // @[OneHot.scala 66:30:@10717.4]
  wire  _T_26504; // @[OneHot.scala 66:30:@10718.4]
  wire  _T_26505; // @[OneHot.scala 66:30:@10719.4]
  wire  _T_26506; // @[OneHot.scala 66:30:@10720.4]
  wire  _T_26507; // @[OneHot.scala 66:30:@10721.4]
  wire  _T_26508; // @[OneHot.scala 66:30:@10722.4]
  wire  _T_26509; // @[OneHot.scala 66:30:@10723.4]
  wire [7:0] _T_26534; // @[Mux.scala 31:69:@10733.4]
  wire [7:0] _T_26535; // @[Mux.scala 31:69:@10734.4]
  wire [7:0] _T_26536; // @[Mux.scala 31:69:@10735.4]
  wire [7:0] _T_26537; // @[Mux.scala 31:69:@10736.4]
  wire [7:0] _T_26538; // @[Mux.scala 31:69:@10737.4]
  wire [7:0] _T_26539; // @[Mux.scala 31:69:@10738.4]
  wire [7:0] _T_26540; // @[Mux.scala 31:69:@10739.4]
  wire [7:0] _T_26541; // @[Mux.scala 31:69:@10740.4]
  wire  _T_26542; // @[OneHot.scala 66:30:@10741.4]
  wire  _T_26543; // @[OneHot.scala 66:30:@10742.4]
  wire  _T_26544; // @[OneHot.scala 66:30:@10743.4]
  wire  _T_26545; // @[OneHot.scala 66:30:@10744.4]
  wire  _T_26546; // @[OneHot.scala 66:30:@10745.4]
  wire  _T_26547; // @[OneHot.scala 66:30:@10746.4]
  wire  _T_26548; // @[OneHot.scala 66:30:@10747.4]
  wire  _T_26549; // @[OneHot.scala 66:30:@10748.4]
  wire [7:0] _T_26590; // @[Mux.scala 19:72:@10764.4]
  wire [7:0] _T_26592; // @[Mux.scala 19:72:@10765.4]
  wire [7:0] _T_26599; // @[Mux.scala 19:72:@10772.4]
  wire [7:0] _T_26601; // @[Mux.scala 19:72:@10773.4]
  wire [7:0] _T_26608; // @[Mux.scala 19:72:@10780.4]
  wire [7:0] _T_26610; // @[Mux.scala 19:72:@10781.4]
  wire [7:0] _T_26617; // @[Mux.scala 19:72:@10788.4]
  wire [7:0] _T_26619; // @[Mux.scala 19:72:@10789.4]
  wire [7:0] _T_26626; // @[Mux.scala 19:72:@10796.4]
  wire [7:0] _T_26628; // @[Mux.scala 19:72:@10797.4]
  wire [7:0] _T_26635; // @[Mux.scala 19:72:@10804.4]
  wire [7:0] _T_26637; // @[Mux.scala 19:72:@10805.4]
  wire [7:0] _T_26644; // @[Mux.scala 19:72:@10812.4]
  wire [7:0] _T_26646; // @[Mux.scala 19:72:@10813.4]
  wire [7:0] _T_26653; // @[Mux.scala 19:72:@10820.4]
  wire [7:0] _T_26655; // @[Mux.scala 19:72:@10821.4]
  wire [7:0] _T_26656; // @[Mux.scala 19:72:@10822.4]
  wire [7:0] _T_26657; // @[Mux.scala 19:72:@10823.4]
  wire [7:0] _T_26658; // @[Mux.scala 19:72:@10824.4]
  wire [7:0] _T_26659; // @[Mux.scala 19:72:@10825.4]
  wire [7:0] _T_26660; // @[Mux.scala 19:72:@10826.4]
  wire [7:0] _T_26661; // @[Mux.scala 19:72:@10827.4]
  wire [7:0] _T_26662; // @[Mux.scala 19:72:@10828.4]
  wire  outputPriorityPorts_0_0; // @[Mux.scala 19:72:@10832.4]
  wire  outputPriorityPorts_0_1; // @[Mux.scala 19:72:@10834.4]
  wire  outputPriorityPorts_0_2; // @[Mux.scala 19:72:@10836.4]
  wire  outputPriorityPorts_0_3; // @[Mux.scala 19:72:@10838.4]
  wire  outputPriorityPorts_0_4; // @[Mux.scala 19:72:@10840.4]
  wire  outputPriorityPorts_0_5; // @[Mux.scala 19:72:@10842.4]
  wire  outputPriorityPorts_0_6; // @[Mux.scala 19:72:@10844.4]
  wire  outputPriorityPorts_0_7; // @[Mux.scala 19:72:@10846.4]
  wire  _T_26742; // @[LoadQueue.scala 298:83:@10857.4]
  wire  _T_26745; // @[LoadQueue.scala 298:83:@10859.4]
  wire  _T_26748; // @[LoadQueue.scala 298:83:@10861.4]
  wire  _T_26751; // @[LoadQueue.scala 298:83:@10863.4]
  wire  _T_26754; // @[LoadQueue.scala 298:83:@10865.4]
  wire  _T_26757; // @[LoadQueue.scala 298:83:@10867.4]
  wire  _T_26760; // @[LoadQueue.scala 298:83:@10869.4]
  wire  _T_26763; // @[LoadQueue.scala 298:83:@10871.4]
  wire [7:0] _T_26814; // @[Mux.scala 31:69:@10901.4]
  wire [7:0] _T_26815; // @[Mux.scala 31:69:@10902.4]
  wire [7:0] _T_26816; // @[Mux.scala 31:69:@10903.4]
  wire [7:0] _T_26817; // @[Mux.scala 31:69:@10904.4]
  wire [7:0] _T_26818; // @[Mux.scala 31:69:@10905.4]
  wire [7:0] _T_26819; // @[Mux.scala 31:69:@10906.4]
  wire [7:0] _T_26820; // @[Mux.scala 31:69:@10907.4]
  wire [7:0] _T_26821; // @[Mux.scala 31:69:@10908.4]
  wire  _T_26822; // @[OneHot.scala 66:30:@10909.4]
  wire  _T_26823; // @[OneHot.scala 66:30:@10910.4]
  wire  _T_26824; // @[OneHot.scala 66:30:@10911.4]
  wire  _T_26825; // @[OneHot.scala 66:30:@10912.4]
  wire  _T_26826; // @[OneHot.scala 66:30:@10913.4]
  wire  _T_26827; // @[OneHot.scala 66:30:@10914.4]
  wire  _T_26828; // @[OneHot.scala 66:30:@10915.4]
  wire  _T_26829; // @[OneHot.scala 66:30:@10916.4]
  wire [7:0] _T_26854; // @[Mux.scala 31:69:@10926.4]
  wire [7:0] _T_26855; // @[Mux.scala 31:69:@10927.4]
  wire [7:0] _T_26856; // @[Mux.scala 31:69:@10928.4]
  wire [7:0] _T_26857; // @[Mux.scala 31:69:@10929.4]
  wire [7:0] _T_26858; // @[Mux.scala 31:69:@10930.4]
  wire [7:0] _T_26859; // @[Mux.scala 31:69:@10931.4]
  wire [7:0] _T_26860; // @[Mux.scala 31:69:@10932.4]
  wire [7:0] _T_26861; // @[Mux.scala 31:69:@10933.4]
  wire  _T_26862; // @[OneHot.scala 66:30:@10934.4]
  wire  _T_26863; // @[OneHot.scala 66:30:@10935.4]
  wire  _T_26864; // @[OneHot.scala 66:30:@10936.4]
  wire  _T_26865; // @[OneHot.scala 66:30:@10937.4]
  wire  _T_26866; // @[OneHot.scala 66:30:@10938.4]
  wire  _T_26867; // @[OneHot.scala 66:30:@10939.4]
  wire  _T_26868; // @[OneHot.scala 66:30:@10940.4]
  wire  _T_26869; // @[OneHot.scala 66:30:@10941.4]
  wire [7:0] _T_26894; // @[Mux.scala 31:69:@10951.4]
  wire [7:0] _T_26895; // @[Mux.scala 31:69:@10952.4]
  wire [7:0] _T_26896; // @[Mux.scala 31:69:@10953.4]
  wire [7:0] _T_26897; // @[Mux.scala 31:69:@10954.4]
  wire [7:0] _T_26898; // @[Mux.scala 31:69:@10955.4]
  wire [7:0] _T_26899; // @[Mux.scala 31:69:@10956.4]
  wire [7:0] _T_26900; // @[Mux.scala 31:69:@10957.4]
  wire [7:0] _T_26901; // @[Mux.scala 31:69:@10958.4]
  wire  _T_26902; // @[OneHot.scala 66:30:@10959.4]
  wire  _T_26903; // @[OneHot.scala 66:30:@10960.4]
  wire  _T_26904; // @[OneHot.scala 66:30:@10961.4]
  wire  _T_26905; // @[OneHot.scala 66:30:@10962.4]
  wire  _T_26906; // @[OneHot.scala 66:30:@10963.4]
  wire  _T_26907; // @[OneHot.scala 66:30:@10964.4]
  wire  _T_26908; // @[OneHot.scala 66:30:@10965.4]
  wire  _T_26909; // @[OneHot.scala 66:30:@10966.4]
  wire [7:0] _T_26934; // @[Mux.scala 31:69:@10976.4]
  wire [7:0] _T_26935; // @[Mux.scala 31:69:@10977.4]
  wire [7:0] _T_26936; // @[Mux.scala 31:69:@10978.4]
  wire [7:0] _T_26937; // @[Mux.scala 31:69:@10979.4]
  wire [7:0] _T_26938; // @[Mux.scala 31:69:@10980.4]
  wire [7:0] _T_26939; // @[Mux.scala 31:69:@10981.4]
  wire [7:0] _T_26940; // @[Mux.scala 31:69:@10982.4]
  wire [7:0] _T_26941; // @[Mux.scala 31:69:@10983.4]
  wire  _T_26942; // @[OneHot.scala 66:30:@10984.4]
  wire  _T_26943; // @[OneHot.scala 66:30:@10985.4]
  wire  _T_26944; // @[OneHot.scala 66:30:@10986.4]
  wire  _T_26945; // @[OneHot.scala 66:30:@10987.4]
  wire  _T_26946; // @[OneHot.scala 66:30:@10988.4]
  wire  _T_26947; // @[OneHot.scala 66:30:@10989.4]
  wire  _T_26948; // @[OneHot.scala 66:30:@10990.4]
  wire  _T_26949; // @[OneHot.scala 66:30:@10991.4]
  wire [7:0] _T_26974; // @[Mux.scala 31:69:@11001.4]
  wire [7:0] _T_26975; // @[Mux.scala 31:69:@11002.4]
  wire [7:0] _T_26976; // @[Mux.scala 31:69:@11003.4]
  wire [7:0] _T_26977; // @[Mux.scala 31:69:@11004.4]
  wire [7:0] _T_26978; // @[Mux.scala 31:69:@11005.4]
  wire [7:0] _T_26979; // @[Mux.scala 31:69:@11006.4]
  wire [7:0] _T_26980; // @[Mux.scala 31:69:@11007.4]
  wire [7:0] _T_26981; // @[Mux.scala 31:69:@11008.4]
  wire  _T_26982; // @[OneHot.scala 66:30:@11009.4]
  wire  _T_26983; // @[OneHot.scala 66:30:@11010.4]
  wire  _T_26984; // @[OneHot.scala 66:30:@11011.4]
  wire  _T_26985; // @[OneHot.scala 66:30:@11012.4]
  wire  _T_26986; // @[OneHot.scala 66:30:@11013.4]
  wire  _T_26987; // @[OneHot.scala 66:30:@11014.4]
  wire  _T_26988; // @[OneHot.scala 66:30:@11015.4]
  wire  _T_26989; // @[OneHot.scala 66:30:@11016.4]
  wire [7:0] _T_27014; // @[Mux.scala 31:69:@11026.4]
  wire [7:0] _T_27015; // @[Mux.scala 31:69:@11027.4]
  wire [7:0] _T_27016; // @[Mux.scala 31:69:@11028.4]
  wire [7:0] _T_27017; // @[Mux.scala 31:69:@11029.4]
  wire [7:0] _T_27018; // @[Mux.scala 31:69:@11030.4]
  wire [7:0] _T_27019; // @[Mux.scala 31:69:@11031.4]
  wire [7:0] _T_27020; // @[Mux.scala 31:69:@11032.4]
  wire [7:0] _T_27021; // @[Mux.scala 31:69:@11033.4]
  wire  _T_27022; // @[OneHot.scala 66:30:@11034.4]
  wire  _T_27023; // @[OneHot.scala 66:30:@11035.4]
  wire  _T_27024; // @[OneHot.scala 66:30:@11036.4]
  wire  _T_27025; // @[OneHot.scala 66:30:@11037.4]
  wire  _T_27026; // @[OneHot.scala 66:30:@11038.4]
  wire  _T_27027; // @[OneHot.scala 66:30:@11039.4]
  wire  _T_27028; // @[OneHot.scala 66:30:@11040.4]
  wire  _T_27029; // @[OneHot.scala 66:30:@11041.4]
  wire [7:0] _T_27054; // @[Mux.scala 31:69:@11051.4]
  wire [7:0] _T_27055; // @[Mux.scala 31:69:@11052.4]
  wire [7:0] _T_27056; // @[Mux.scala 31:69:@11053.4]
  wire [7:0] _T_27057; // @[Mux.scala 31:69:@11054.4]
  wire [7:0] _T_27058; // @[Mux.scala 31:69:@11055.4]
  wire [7:0] _T_27059; // @[Mux.scala 31:69:@11056.4]
  wire [7:0] _T_27060; // @[Mux.scala 31:69:@11057.4]
  wire [7:0] _T_27061; // @[Mux.scala 31:69:@11058.4]
  wire  _T_27062; // @[OneHot.scala 66:30:@11059.4]
  wire  _T_27063; // @[OneHot.scala 66:30:@11060.4]
  wire  _T_27064; // @[OneHot.scala 66:30:@11061.4]
  wire  _T_27065; // @[OneHot.scala 66:30:@11062.4]
  wire  _T_27066; // @[OneHot.scala 66:30:@11063.4]
  wire  _T_27067; // @[OneHot.scala 66:30:@11064.4]
  wire  _T_27068; // @[OneHot.scala 66:30:@11065.4]
  wire  _T_27069; // @[OneHot.scala 66:30:@11066.4]
  wire [7:0] _T_27094; // @[Mux.scala 31:69:@11076.4]
  wire [7:0] _T_27095; // @[Mux.scala 31:69:@11077.4]
  wire [7:0] _T_27096; // @[Mux.scala 31:69:@11078.4]
  wire [7:0] _T_27097; // @[Mux.scala 31:69:@11079.4]
  wire [7:0] _T_27098; // @[Mux.scala 31:69:@11080.4]
  wire [7:0] _T_27099; // @[Mux.scala 31:69:@11081.4]
  wire [7:0] _T_27100; // @[Mux.scala 31:69:@11082.4]
  wire [7:0] _T_27101; // @[Mux.scala 31:69:@11083.4]
  wire  _T_27102; // @[OneHot.scala 66:30:@11084.4]
  wire  _T_27103; // @[OneHot.scala 66:30:@11085.4]
  wire  _T_27104; // @[OneHot.scala 66:30:@11086.4]
  wire  _T_27105; // @[OneHot.scala 66:30:@11087.4]
  wire  _T_27106; // @[OneHot.scala 66:30:@11088.4]
  wire  _T_27107; // @[OneHot.scala 66:30:@11089.4]
  wire  _T_27108; // @[OneHot.scala 66:30:@11090.4]
  wire  _T_27109; // @[OneHot.scala 66:30:@11091.4]
  wire [7:0] _T_27150; // @[Mux.scala 19:72:@11107.4]
  wire [7:0] _T_27152; // @[Mux.scala 19:72:@11108.4]
  wire [7:0] _T_27159; // @[Mux.scala 19:72:@11115.4]
  wire [7:0] _T_27161; // @[Mux.scala 19:72:@11116.4]
  wire [7:0] _T_27168; // @[Mux.scala 19:72:@11123.4]
  wire [7:0] _T_27170; // @[Mux.scala 19:72:@11124.4]
  wire [7:0] _T_27177; // @[Mux.scala 19:72:@11131.4]
  wire [7:0] _T_27179; // @[Mux.scala 19:72:@11132.4]
  wire [7:0] _T_27186; // @[Mux.scala 19:72:@11139.4]
  wire [7:0] _T_27188; // @[Mux.scala 19:72:@11140.4]
  wire [7:0] _T_27195; // @[Mux.scala 19:72:@11147.4]
  wire [7:0] _T_27197; // @[Mux.scala 19:72:@11148.4]
  wire [7:0] _T_27204; // @[Mux.scala 19:72:@11155.4]
  wire [7:0] _T_27206; // @[Mux.scala 19:72:@11156.4]
  wire [7:0] _T_27213; // @[Mux.scala 19:72:@11163.4]
  wire [7:0] _T_27215; // @[Mux.scala 19:72:@11164.4]
  wire [7:0] _T_27216; // @[Mux.scala 19:72:@11165.4]
  wire [7:0] _T_27217; // @[Mux.scala 19:72:@11166.4]
  wire [7:0] _T_27218; // @[Mux.scala 19:72:@11167.4]
  wire [7:0] _T_27219; // @[Mux.scala 19:72:@11168.4]
  wire [7:0] _T_27220; // @[Mux.scala 19:72:@11169.4]
  wire [7:0] _T_27221; // @[Mux.scala 19:72:@11170.4]
  wire [7:0] _T_27222; // @[Mux.scala 19:72:@11171.4]
  wire  inputPriorityPorts_1_0; // @[Mux.scala 19:72:@11175.4]
  wire  inputPriorityPorts_1_1; // @[Mux.scala 19:72:@11177.4]
  wire  inputPriorityPorts_1_2; // @[Mux.scala 19:72:@11179.4]
  wire  inputPriorityPorts_1_3; // @[Mux.scala 19:72:@11181.4]
  wire  inputPriorityPorts_1_4; // @[Mux.scala 19:72:@11183.4]
  wire  inputPriorityPorts_1_5; // @[Mux.scala 19:72:@11185.4]
  wire  inputPriorityPorts_1_6; // @[Mux.scala 19:72:@11187.4]
  wire  inputPriorityPorts_1_7; // @[Mux.scala 19:72:@11189.4]
  wire [7:0] _T_27336; // @[Mux.scala 31:69:@11219.4]
  wire [7:0] _T_27337; // @[Mux.scala 31:69:@11220.4]
  wire [7:0] _T_27338; // @[Mux.scala 31:69:@11221.4]
  wire [7:0] _T_27339; // @[Mux.scala 31:69:@11222.4]
  wire [7:0] _T_27340; // @[Mux.scala 31:69:@11223.4]
  wire [7:0] _T_27341; // @[Mux.scala 31:69:@11224.4]
  wire [7:0] _T_27342; // @[Mux.scala 31:69:@11225.4]
  wire [7:0] _T_27343; // @[Mux.scala 31:69:@11226.4]
  wire  _T_27344; // @[OneHot.scala 66:30:@11227.4]
  wire  _T_27345; // @[OneHot.scala 66:30:@11228.4]
  wire  _T_27346; // @[OneHot.scala 66:30:@11229.4]
  wire  _T_27347; // @[OneHot.scala 66:30:@11230.4]
  wire  _T_27348; // @[OneHot.scala 66:30:@11231.4]
  wire  _T_27349; // @[OneHot.scala 66:30:@11232.4]
  wire  _T_27350; // @[OneHot.scala 66:30:@11233.4]
  wire  _T_27351; // @[OneHot.scala 66:30:@11234.4]
  wire [7:0] _T_27376; // @[Mux.scala 31:69:@11244.4]
  wire [7:0] _T_27377; // @[Mux.scala 31:69:@11245.4]
  wire [7:0] _T_27378; // @[Mux.scala 31:69:@11246.4]
  wire [7:0] _T_27379; // @[Mux.scala 31:69:@11247.4]
  wire [7:0] _T_27380; // @[Mux.scala 31:69:@11248.4]
  wire [7:0] _T_27381; // @[Mux.scala 31:69:@11249.4]
  wire [7:0] _T_27382; // @[Mux.scala 31:69:@11250.4]
  wire [7:0] _T_27383; // @[Mux.scala 31:69:@11251.4]
  wire  _T_27384; // @[OneHot.scala 66:30:@11252.4]
  wire  _T_27385; // @[OneHot.scala 66:30:@11253.4]
  wire  _T_27386; // @[OneHot.scala 66:30:@11254.4]
  wire  _T_27387; // @[OneHot.scala 66:30:@11255.4]
  wire  _T_27388; // @[OneHot.scala 66:30:@11256.4]
  wire  _T_27389; // @[OneHot.scala 66:30:@11257.4]
  wire  _T_27390; // @[OneHot.scala 66:30:@11258.4]
  wire  _T_27391; // @[OneHot.scala 66:30:@11259.4]
  wire [7:0] _T_27416; // @[Mux.scala 31:69:@11269.4]
  wire [7:0] _T_27417; // @[Mux.scala 31:69:@11270.4]
  wire [7:0] _T_27418; // @[Mux.scala 31:69:@11271.4]
  wire [7:0] _T_27419; // @[Mux.scala 31:69:@11272.4]
  wire [7:0] _T_27420; // @[Mux.scala 31:69:@11273.4]
  wire [7:0] _T_27421; // @[Mux.scala 31:69:@11274.4]
  wire [7:0] _T_27422; // @[Mux.scala 31:69:@11275.4]
  wire [7:0] _T_27423; // @[Mux.scala 31:69:@11276.4]
  wire  _T_27424; // @[OneHot.scala 66:30:@11277.4]
  wire  _T_27425; // @[OneHot.scala 66:30:@11278.4]
  wire  _T_27426; // @[OneHot.scala 66:30:@11279.4]
  wire  _T_27427; // @[OneHot.scala 66:30:@11280.4]
  wire  _T_27428; // @[OneHot.scala 66:30:@11281.4]
  wire  _T_27429; // @[OneHot.scala 66:30:@11282.4]
  wire  _T_27430; // @[OneHot.scala 66:30:@11283.4]
  wire  _T_27431; // @[OneHot.scala 66:30:@11284.4]
  wire [7:0] _T_27456; // @[Mux.scala 31:69:@11294.4]
  wire [7:0] _T_27457; // @[Mux.scala 31:69:@11295.4]
  wire [7:0] _T_27458; // @[Mux.scala 31:69:@11296.4]
  wire [7:0] _T_27459; // @[Mux.scala 31:69:@11297.4]
  wire [7:0] _T_27460; // @[Mux.scala 31:69:@11298.4]
  wire [7:0] _T_27461; // @[Mux.scala 31:69:@11299.4]
  wire [7:0] _T_27462; // @[Mux.scala 31:69:@11300.4]
  wire [7:0] _T_27463; // @[Mux.scala 31:69:@11301.4]
  wire  _T_27464; // @[OneHot.scala 66:30:@11302.4]
  wire  _T_27465; // @[OneHot.scala 66:30:@11303.4]
  wire  _T_27466; // @[OneHot.scala 66:30:@11304.4]
  wire  _T_27467; // @[OneHot.scala 66:30:@11305.4]
  wire  _T_27468; // @[OneHot.scala 66:30:@11306.4]
  wire  _T_27469; // @[OneHot.scala 66:30:@11307.4]
  wire  _T_27470; // @[OneHot.scala 66:30:@11308.4]
  wire  _T_27471; // @[OneHot.scala 66:30:@11309.4]
  wire [7:0] _T_27496; // @[Mux.scala 31:69:@11319.4]
  wire [7:0] _T_27497; // @[Mux.scala 31:69:@11320.4]
  wire [7:0] _T_27498; // @[Mux.scala 31:69:@11321.4]
  wire [7:0] _T_27499; // @[Mux.scala 31:69:@11322.4]
  wire [7:0] _T_27500; // @[Mux.scala 31:69:@11323.4]
  wire [7:0] _T_27501; // @[Mux.scala 31:69:@11324.4]
  wire [7:0] _T_27502; // @[Mux.scala 31:69:@11325.4]
  wire [7:0] _T_27503; // @[Mux.scala 31:69:@11326.4]
  wire  _T_27504; // @[OneHot.scala 66:30:@11327.4]
  wire  _T_27505; // @[OneHot.scala 66:30:@11328.4]
  wire  _T_27506; // @[OneHot.scala 66:30:@11329.4]
  wire  _T_27507; // @[OneHot.scala 66:30:@11330.4]
  wire  _T_27508; // @[OneHot.scala 66:30:@11331.4]
  wire  _T_27509; // @[OneHot.scala 66:30:@11332.4]
  wire  _T_27510; // @[OneHot.scala 66:30:@11333.4]
  wire  _T_27511; // @[OneHot.scala 66:30:@11334.4]
  wire [7:0] _T_27536; // @[Mux.scala 31:69:@11344.4]
  wire [7:0] _T_27537; // @[Mux.scala 31:69:@11345.4]
  wire [7:0] _T_27538; // @[Mux.scala 31:69:@11346.4]
  wire [7:0] _T_27539; // @[Mux.scala 31:69:@11347.4]
  wire [7:0] _T_27540; // @[Mux.scala 31:69:@11348.4]
  wire [7:0] _T_27541; // @[Mux.scala 31:69:@11349.4]
  wire [7:0] _T_27542; // @[Mux.scala 31:69:@11350.4]
  wire [7:0] _T_27543; // @[Mux.scala 31:69:@11351.4]
  wire  _T_27544; // @[OneHot.scala 66:30:@11352.4]
  wire  _T_27545; // @[OneHot.scala 66:30:@11353.4]
  wire  _T_27546; // @[OneHot.scala 66:30:@11354.4]
  wire  _T_27547; // @[OneHot.scala 66:30:@11355.4]
  wire  _T_27548; // @[OneHot.scala 66:30:@11356.4]
  wire  _T_27549; // @[OneHot.scala 66:30:@11357.4]
  wire  _T_27550; // @[OneHot.scala 66:30:@11358.4]
  wire  _T_27551; // @[OneHot.scala 66:30:@11359.4]
  wire [7:0] _T_27576; // @[Mux.scala 31:69:@11369.4]
  wire [7:0] _T_27577; // @[Mux.scala 31:69:@11370.4]
  wire [7:0] _T_27578; // @[Mux.scala 31:69:@11371.4]
  wire [7:0] _T_27579; // @[Mux.scala 31:69:@11372.4]
  wire [7:0] _T_27580; // @[Mux.scala 31:69:@11373.4]
  wire [7:0] _T_27581; // @[Mux.scala 31:69:@11374.4]
  wire [7:0] _T_27582; // @[Mux.scala 31:69:@11375.4]
  wire [7:0] _T_27583; // @[Mux.scala 31:69:@11376.4]
  wire  _T_27584; // @[OneHot.scala 66:30:@11377.4]
  wire  _T_27585; // @[OneHot.scala 66:30:@11378.4]
  wire  _T_27586; // @[OneHot.scala 66:30:@11379.4]
  wire  _T_27587; // @[OneHot.scala 66:30:@11380.4]
  wire  _T_27588; // @[OneHot.scala 66:30:@11381.4]
  wire  _T_27589; // @[OneHot.scala 66:30:@11382.4]
  wire  _T_27590; // @[OneHot.scala 66:30:@11383.4]
  wire  _T_27591; // @[OneHot.scala 66:30:@11384.4]
  wire [7:0] _T_27616; // @[Mux.scala 31:69:@11394.4]
  wire [7:0] _T_27617; // @[Mux.scala 31:69:@11395.4]
  wire [7:0] _T_27618; // @[Mux.scala 31:69:@11396.4]
  wire [7:0] _T_27619; // @[Mux.scala 31:69:@11397.4]
  wire [7:0] _T_27620; // @[Mux.scala 31:69:@11398.4]
  wire [7:0] _T_27621; // @[Mux.scala 31:69:@11399.4]
  wire [7:0] _T_27622; // @[Mux.scala 31:69:@11400.4]
  wire [7:0] _T_27623; // @[Mux.scala 31:69:@11401.4]
  wire  _T_27624; // @[OneHot.scala 66:30:@11402.4]
  wire  _T_27625; // @[OneHot.scala 66:30:@11403.4]
  wire  _T_27626; // @[OneHot.scala 66:30:@11404.4]
  wire  _T_27627; // @[OneHot.scala 66:30:@11405.4]
  wire  _T_27628; // @[OneHot.scala 66:30:@11406.4]
  wire  _T_27629; // @[OneHot.scala 66:30:@11407.4]
  wire  _T_27630; // @[OneHot.scala 66:30:@11408.4]
  wire  _T_27631; // @[OneHot.scala 66:30:@11409.4]
  wire [7:0] _T_27672; // @[Mux.scala 19:72:@11425.4]
  wire [7:0] _T_27674; // @[Mux.scala 19:72:@11426.4]
  wire [7:0] _T_27681; // @[Mux.scala 19:72:@11433.4]
  wire [7:0] _T_27683; // @[Mux.scala 19:72:@11434.4]
  wire [7:0] _T_27690; // @[Mux.scala 19:72:@11441.4]
  wire [7:0] _T_27692; // @[Mux.scala 19:72:@11442.4]
  wire [7:0] _T_27699; // @[Mux.scala 19:72:@11449.4]
  wire [7:0] _T_27701; // @[Mux.scala 19:72:@11450.4]
  wire [7:0] _T_27708; // @[Mux.scala 19:72:@11457.4]
  wire [7:0] _T_27710; // @[Mux.scala 19:72:@11458.4]
  wire [7:0] _T_27717; // @[Mux.scala 19:72:@11465.4]
  wire [7:0] _T_27719; // @[Mux.scala 19:72:@11466.4]
  wire [7:0] _T_27726; // @[Mux.scala 19:72:@11473.4]
  wire [7:0] _T_27728; // @[Mux.scala 19:72:@11474.4]
  wire [7:0] _T_27735; // @[Mux.scala 19:72:@11481.4]
  wire [7:0] _T_27737; // @[Mux.scala 19:72:@11482.4]
  wire [7:0] _T_27738; // @[Mux.scala 19:72:@11483.4]
  wire [7:0] _T_27739; // @[Mux.scala 19:72:@11484.4]
  wire [7:0] _T_27740; // @[Mux.scala 19:72:@11485.4]
  wire [7:0] _T_27741; // @[Mux.scala 19:72:@11486.4]
  wire [7:0] _T_27742; // @[Mux.scala 19:72:@11487.4]
  wire [7:0] _T_27743; // @[Mux.scala 19:72:@11488.4]
  wire [7:0] _T_27744; // @[Mux.scala 19:72:@11489.4]
  wire  outputPriorityPorts_1_0; // @[Mux.scala 19:72:@11493.4]
  wire  outputPriorityPorts_1_1; // @[Mux.scala 19:72:@11495.4]
  wire  outputPriorityPorts_1_2; // @[Mux.scala 19:72:@11497.4]
  wire  outputPriorityPorts_1_3; // @[Mux.scala 19:72:@11499.4]
  wire  outputPriorityPorts_1_4; // @[Mux.scala 19:72:@11501.4]
  wire  outputPriorityPorts_1_5; // @[Mux.scala 19:72:@11503.4]
  wire  outputPriorityPorts_1_6; // @[Mux.scala 19:72:@11505.4]
  wire  outputPriorityPorts_1_7; // @[Mux.scala 19:72:@11507.4]
  wire  _T_27823; // @[LoadQueue.scala 313:47:@11521.6]
  wire  _T_27824; // @[LoadQueue.scala 313:47:@11522.6]
  wire  _T_27835; // @[LoadQueue.scala 314:26:@11527.6]
  wire [1:0] _T_27836; // @[OneHot.scala 18:45:@11529.8]
  wire  _T_27837; // @[CircuitMath.scala 30:8:@11530.8]
  wire [31:0] _GEN_611; // @[LoadQueue.scala 315:29:@11531.8]
  wire [31:0] _GEN_612; // @[LoadQueue.scala 314:36:@11528.6]
  wire  _GEN_613; // @[LoadQueue.scala 314:36:@11528.6]
  wire  _GEN_614; // @[LoadQueue.scala 308:34:@11517.4]
  wire [31:0] _GEN_615; // @[LoadQueue.scala 308:34:@11517.4]
  wire  _T_27841; // @[LoadQueue.scala 313:47:@11539.6]
  wire  _T_27842; // @[LoadQueue.scala 313:47:@11540.6]
  wire  _T_27853; // @[LoadQueue.scala 314:26:@11545.6]
  wire [1:0] _T_27854; // @[OneHot.scala 18:45:@11547.8]
  wire  _T_27855; // @[CircuitMath.scala 30:8:@11548.8]
  wire [31:0] _GEN_617; // @[LoadQueue.scala 315:29:@11549.8]
  wire [31:0] _GEN_618; // @[LoadQueue.scala 314:36:@11546.6]
  wire  _GEN_619; // @[LoadQueue.scala 314:36:@11546.6]
  wire  _GEN_620; // @[LoadQueue.scala 308:34:@11535.4]
  wire [31:0] _GEN_621; // @[LoadQueue.scala 308:34:@11535.4]
  wire  _T_27859; // @[LoadQueue.scala 313:47:@11557.6]
  wire  _T_27860; // @[LoadQueue.scala 313:47:@11558.6]
  wire  _T_27871; // @[LoadQueue.scala 314:26:@11563.6]
  wire [1:0] _T_27872; // @[OneHot.scala 18:45:@11565.8]
  wire  _T_27873; // @[CircuitMath.scala 30:8:@11566.8]
  wire [31:0] _GEN_623; // @[LoadQueue.scala 315:29:@11567.8]
  wire [31:0] _GEN_624; // @[LoadQueue.scala 314:36:@11564.6]
  wire  _GEN_625; // @[LoadQueue.scala 314:36:@11564.6]
  wire  _GEN_626; // @[LoadQueue.scala 308:34:@11553.4]
  wire [31:0] _GEN_627; // @[LoadQueue.scala 308:34:@11553.4]
  wire  _T_27877; // @[LoadQueue.scala 313:47:@11575.6]
  wire  _T_27878; // @[LoadQueue.scala 313:47:@11576.6]
  wire  _T_27889; // @[LoadQueue.scala 314:26:@11581.6]
  wire [1:0] _T_27890; // @[OneHot.scala 18:45:@11583.8]
  wire  _T_27891; // @[CircuitMath.scala 30:8:@11584.8]
  wire [31:0] _GEN_629; // @[LoadQueue.scala 315:29:@11585.8]
  wire [31:0] _GEN_630; // @[LoadQueue.scala 314:36:@11582.6]
  wire  _GEN_631; // @[LoadQueue.scala 314:36:@11582.6]
  wire  _GEN_632; // @[LoadQueue.scala 308:34:@11571.4]
  wire [31:0] _GEN_633; // @[LoadQueue.scala 308:34:@11571.4]
  wire  _T_27895; // @[LoadQueue.scala 313:47:@11593.6]
  wire  _T_27896; // @[LoadQueue.scala 313:47:@11594.6]
  wire  _T_27907; // @[LoadQueue.scala 314:26:@11599.6]
  wire [1:0] _T_27908; // @[OneHot.scala 18:45:@11601.8]
  wire  _T_27909; // @[CircuitMath.scala 30:8:@11602.8]
  wire [31:0] _GEN_635; // @[LoadQueue.scala 315:29:@11603.8]
  wire [31:0] _GEN_636; // @[LoadQueue.scala 314:36:@11600.6]
  wire  _GEN_637; // @[LoadQueue.scala 314:36:@11600.6]
  wire  _GEN_638; // @[LoadQueue.scala 308:34:@11589.4]
  wire [31:0] _GEN_639; // @[LoadQueue.scala 308:34:@11589.4]
  wire  _T_27913; // @[LoadQueue.scala 313:47:@11611.6]
  wire  _T_27914; // @[LoadQueue.scala 313:47:@11612.6]
  wire  _T_27925; // @[LoadQueue.scala 314:26:@11617.6]
  wire [1:0] _T_27926; // @[OneHot.scala 18:45:@11619.8]
  wire  _T_27927; // @[CircuitMath.scala 30:8:@11620.8]
  wire [31:0] _GEN_641; // @[LoadQueue.scala 315:29:@11621.8]
  wire [31:0] _GEN_642; // @[LoadQueue.scala 314:36:@11618.6]
  wire  _GEN_643; // @[LoadQueue.scala 314:36:@11618.6]
  wire  _GEN_644; // @[LoadQueue.scala 308:34:@11607.4]
  wire [31:0] _GEN_645; // @[LoadQueue.scala 308:34:@11607.4]
  wire  _T_27931; // @[LoadQueue.scala 313:47:@11629.6]
  wire  _T_27932; // @[LoadQueue.scala 313:47:@11630.6]
  wire  _T_27943; // @[LoadQueue.scala 314:26:@11635.6]
  wire [1:0] _T_27944; // @[OneHot.scala 18:45:@11637.8]
  wire  _T_27945; // @[CircuitMath.scala 30:8:@11638.8]
  wire [31:0] _GEN_647; // @[LoadQueue.scala 315:29:@11639.8]
  wire [31:0] _GEN_648; // @[LoadQueue.scala 314:36:@11636.6]
  wire  _GEN_649; // @[LoadQueue.scala 314:36:@11636.6]
  wire  _GEN_650; // @[LoadQueue.scala 308:34:@11625.4]
  wire [31:0] _GEN_651; // @[LoadQueue.scala 308:34:@11625.4]
  wire  _T_27949; // @[LoadQueue.scala 313:47:@11647.6]
  wire  _T_27950; // @[LoadQueue.scala 313:47:@11648.6]
  wire  _T_27961; // @[LoadQueue.scala 314:26:@11653.6]
  wire [1:0] _T_27962; // @[OneHot.scala 18:45:@11655.8]
  wire  _T_27963; // @[CircuitMath.scala 30:8:@11656.8]
  wire [31:0] _GEN_653; // @[LoadQueue.scala 315:29:@11657.8]
  wire [31:0] _GEN_654; // @[LoadQueue.scala 314:36:@11654.6]
  wire  _GEN_655; // @[LoadQueue.scala 314:36:@11654.6]
  wire  _GEN_656; // @[LoadQueue.scala 308:34:@11643.4]
  wire [31:0] _GEN_657; // @[LoadQueue.scala 308:34:@11643.4]
  wire  _T_27979; // @[LoadQueue.scala 326:108:@11662.4]
  wire  _T_27981; // @[LoadQueue.scala 327:34:@11663.4]
  wire  _T_27982; // @[LoadQueue.scala 327:31:@11664.4]
  wire  _T_27983; // @[LoadQueue.scala 327:63:@11665.4]
  wire  _T_27984; // @[LoadQueue.scala 326:108:@11666.4]
  wire  _T_27987; // @[LoadQueue.scala 327:31:@11668.4]
  wire  _T_27988; // @[LoadQueue.scala 327:63:@11669.4]
  wire  loadCompleting_0; // @[LoadQueue.scala 328:51:@11674.4]
  wire  _T_28000; // @[LoadQueue.scala 326:108:@11676.4]
  wire  _T_28002; // @[LoadQueue.scala 327:34:@11677.4]
  wire  _T_28003; // @[LoadQueue.scala 327:31:@11678.4]
  wire  _T_28004; // @[LoadQueue.scala 327:63:@11679.4]
  wire  _T_28005; // @[LoadQueue.scala 326:108:@11680.4]
  wire  _T_28008; // @[LoadQueue.scala 327:31:@11682.4]
  wire  _T_28009; // @[LoadQueue.scala 327:63:@11683.4]
  wire  loadCompleting_1; // @[LoadQueue.scala 328:51:@11688.4]
  wire  _T_28021; // @[LoadQueue.scala 326:108:@11690.4]
  wire  _T_28023; // @[LoadQueue.scala 327:34:@11691.4]
  wire  _T_28024; // @[LoadQueue.scala 327:31:@11692.4]
  wire  _T_28025; // @[LoadQueue.scala 327:63:@11693.4]
  wire  _T_28026; // @[LoadQueue.scala 326:108:@11694.4]
  wire  _T_28029; // @[LoadQueue.scala 327:31:@11696.4]
  wire  _T_28030; // @[LoadQueue.scala 327:63:@11697.4]
  wire  loadCompleting_2; // @[LoadQueue.scala 328:51:@11702.4]
  wire  _T_28042; // @[LoadQueue.scala 326:108:@11704.4]
  wire  _T_28044; // @[LoadQueue.scala 327:34:@11705.4]
  wire  _T_28045; // @[LoadQueue.scala 327:31:@11706.4]
  wire  _T_28046; // @[LoadQueue.scala 327:63:@11707.4]
  wire  _T_28047; // @[LoadQueue.scala 326:108:@11708.4]
  wire  _T_28050; // @[LoadQueue.scala 327:31:@11710.4]
  wire  _T_28051; // @[LoadQueue.scala 327:63:@11711.4]
  wire  loadCompleting_3; // @[LoadQueue.scala 328:51:@11716.4]
  wire  _T_28063; // @[LoadQueue.scala 326:108:@11718.4]
  wire  _T_28065; // @[LoadQueue.scala 327:34:@11719.4]
  wire  _T_28066; // @[LoadQueue.scala 327:31:@11720.4]
  wire  _T_28067; // @[LoadQueue.scala 327:63:@11721.4]
  wire  _T_28068; // @[LoadQueue.scala 326:108:@11722.4]
  wire  _T_28071; // @[LoadQueue.scala 327:31:@11724.4]
  wire  _T_28072; // @[LoadQueue.scala 327:63:@11725.4]
  wire  loadCompleting_4; // @[LoadQueue.scala 328:51:@11730.4]
  wire  _T_28084; // @[LoadQueue.scala 326:108:@11732.4]
  wire  _T_28086; // @[LoadQueue.scala 327:34:@11733.4]
  wire  _T_28087; // @[LoadQueue.scala 327:31:@11734.4]
  wire  _T_28088; // @[LoadQueue.scala 327:63:@11735.4]
  wire  _T_28089; // @[LoadQueue.scala 326:108:@11736.4]
  wire  _T_28092; // @[LoadQueue.scala 327:31:@11738.4]
  wire  _T_28093; // @[LoadQueue.scala 327:63:@11739.4]
  wire  loadCompleting_5; // @[LoadQueue.scala 328:51:@11744.4]
  wire  _T_28105; // @[LoadQueue.scala 326:108:@11746.4]
  wire  _T_28107; // @[LoadQueue.scala 327:34:@11747.4]
  wire  _T_28108; // @[LoadQueue.scala 327:31:@11748.4]
  wire  _T_28109; // @[LoadQueue.scala 327:63:@11749.4]
  wire  _T_28110; // @[LoadQueue.scala 326:108:@11750.4]
  wire  _T_28113; // @[LoadQueue.scala 327:31:@11752.4]
  wire  _T_28114; // @[LoadQueue.scala 327:63:@11753.4]
  wire  loadCompleting_6; // @[LoadQueue.scala 328:51:@11758.4]
  wire  _T_28126; // @[LoadQueue.scala 326:108:@11760.4]
  wire  _T_28128; // @[LoadQueue.scala 327:34:@11761.4]
  wire  _T_28129; // @[LoadQueue.scala 327:31:@11762.4]
  wire  _T_28130; // @[LoadQueue.scala 327:63:@11763.4]
  wire  _T_28131; // @[LoadQueue.scala 326:108:@11764.4]
  wire  _T_28134; // @[LoadQueue.scala 327:31:@11766.4]
  wire  _T_28135; // @[LoadQueue.scala 327:63:@11767.4]
  wire  loadCompleting_7; // @[LoadQueue.scala 328:51:@11772.4]
  wire  _GEN_658; // @[LoadQueue.scala 337:46:@11778.6]
  wire  _GEN_659; // @[LoadQueue.scala 335:34:@11774.4]
  wire  _GEN_660; // @[LoadQueue.scala 337:46:@11785.6]
  wire  _GEN_661; // @[LoadQueue.scala 335:34:@11781.4]
  wire  _GEN_662; // @[LoadQueue.scala 337:46:@11792.6]
  wire  _GEN_663; // @[LoadQueue.scala 335:34:@11788.4]
  wire  _GEN_664; // @[LoadQueue.scala 337:46:@11799.6]
  wire  _GEN_665; // @[LoadQueue.scala 335:34:@11795.4]
  wire  _GEN_666; // @[LoadQueue.scala 337:46:@11806.6]
  wire  _GEN_667; // @[LoadQueue.scala 335:34:@11802.4]
  wire  _GEN_668; // @[LoadQueue.scala 337:46:@11813.6]
  wire  _GEN_669; // @[LoadQueue.scala 335:34:@11809.4]
  wire  _GEN_670; // @[LoadQueue.scala 337:46:@11820.6]
  wire  _GEN_671; // @[LoadQueue.scala 335:34:@11816.4]
  wire  _GEN_672; // @[LoadQueue.scala 337:46:@11827.6]
  wire  _GEN_673; // @[LoadQueue.scala 335:34:@11823.4]
  wire  _T_28211; // @[LoadQueue.scala 348:24:@11864.4]
  wire  _T_28212; // @[LoadQueue.scala 348:24:@11865.4]
  wire  _T_28213; // @[LoadQueue.scala 348:24:@11866.4]
  wire  _T_28214; // @[LoadQueue.scala 348:24:@11867.4]
  wire  _T_28215; // @[LoadQueue.scala 348:24:@11868.4]
  wire  _T_28216; // @[LoadQueue.scala 348:24:@11869.4]
  wire  _T_28217; // @[LoadQueue.scala 348:24:@11870.4]
  wire [2:0] _T_28226; // @[Mux.scala 31:69:@11872.6]
  wire [2:0] _T_28227; // @[Mux.scala 31:69:@11873.6]
  wire [2:0] _T_28228; // @[Mux.scala 31:69:@11874.6]
  wire [2:0] _T_28229; // @[Mux.scala 31:69:@11875.6]
  wire [2:0] _T_28230; // @[Mux.scala 31:69:@11876.6]
  wire [2:0] _T_28231; // @[Mux.scala 31:69:@11877.6]
  wire [2:0] _T_28232; // @[Mux.scala 31:69:@11878.6]
  wire [31:0] _GEN_675; // @[LoadQueue.scala 349:37:@11879.6]
  wire [31:0] _GEN_676; // @[LoadQueue.scala 349:37:@11879.6]
  wire [31:0] _GEN_677; // @[LoadQueue.scala 349:37:@11879.6]
  wire [31:0] _GEN_678; // @[LoadQueue.scala 349:37:@11879.6]
  wire [31:0] _GEN_679; // @[LoadQueue.scala 349:37:@11879.6]
  wire [31:0] _GEN_680; // @[LoadQueue.scala 349:37:@11879.6]
  wire [31:0] _GEN_681; // @[LoadQueue.scala 349:37:@11879.6]
  wire  _T_28287; // @[LoadQueue.scala 348:24:@11920.4]
  wire  _T_28288; // @[LoadQueue.scala 348:24:@11921.4]
  wire  _T_28289; // @[LoadQueue.scala 348:24:@11922.4]
  wire  _T_28290; // @[LoadQueue.scala 348:24:@11923.4]
  wire  _T_28291; // @[LoadQueue.scala 348:24:@11924.4]
  wire  _T_28292; // @[LoadQueue.scala 348:24:@11925.4]
  wire  _T_28293; // @[LoadQueue.scala 348:24:@11926.4]
  wire [2:0] _T_28302; // @[Mux.scala 31:69:@11928.6]
  wire [2:0] _T_28303; // @[Mux.scala 31:69:@11929.6]
  wire [2:0] _T_28304; // @[Mux.scala 31:69:@11930.6]
  wire [2:0] _T_28305; // @[Mux.scala 31:69:@11931.6]
  wire [2:0] _T_28306; // @[Mux.scala 31:69:@11932.6]
  wire [2:0] _T_28307; // @[Mux.scala 31:69:@11933.6]
  wire [2:0] _T_28308; // @[Mux.scala 31:69:@11934.6]
  wire [31:0] _GEN_685; // @[LoadQueue.scala 349:37:@11935.6]
  wire [31:0] _GEN_686; // @[LoadQueue.scala 349:37:@11935.6]
  wire [31:0] _GEN_687; // @[LoadQueue.scala 349:37:@11935.6]
  wire [31:0] _GEN_688; // @[LoadQueue.scala 349:37:@11935.6]
  wire [31:0] _GEN_689; // @[LoadQueue.scala 349:37:@11935.6]
  wire [31:0] _GEN_690; // @[LoadQueue.scala 349:37:@11935.6]
  wire [31:0] _GEN_691; // @[LoadQueue.scala 349:37:@11935.6]
  wire  _GEN_695; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_696; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_697; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_698; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_699; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_700; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_701; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_703; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_704; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_705; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_706; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_707; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_708; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _GEN_709; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _T_28319; // @[LoadQueue.scala 363:29:@11942.4]
  wire  _T_28320; // @[LoadQueue.scala 363:63:@11943.4]
  wire  _T_28322; // @[LoadQueue.scala 363:75:@11944.4]
  wire  _T_28323; // @[LoadQueue.scala 363:72:@11945.4]
  wire  _T_28324; // @[LoadQueue.scala 363:54:@11946.4]
  wire [3:0] _T_28327; // @[util.scala 10:8:@11948.6]
  wire [3:0] _GEN_144; // @[util.scala 10:14:@11949.6]
  wire [3:0] _T_28328; // @[util.scala 10:14:@11949.6]
  wire [3:0] _GEN_710; // @[LoadQueue.scala 363:91:@11947.4]
  wire [2:0] _GEN_760; // @[util.scala 10:8:@11953.6]
  wire [3:0] _T_28330; // @[util.scala 10:8:@11953.6]
  wire [3:0] _GEN_145; // @[util.scala 10:14:@11954.6]
  wire [3:0] _T_28331; // @[util.scala 10:14:@11954.6]
  wire [3:0] _GEN_711; // @[LoadQueue.scala 367:20:@11952.4]
  wire  _T_28333; // @[LoadQueue.scala 371:82:@11957.4]
  wire  _T_28334; // @[LoadQueue.scala 371:79:@11958.4]
  wire  _T_28336; // @[LoadQueue.scala 371:82:@11959.4]
  wire  _T_28337; // @[LoadQueue.scala 371:79:@11960.4]
  wire  _T_28339; // @[LoadQueue.scala 371:82:@11961.4]
  wire  _T_28340; // @[LoadQueue.scala 371:79:@11962.4]
  wire  _T_28342; // @[LoadQueue.scala 371:82:@11963.4]
  wire  _T_28343; // @[LoadQueue.scala 371:79:@11964.4]
  wire  _T_28345; // @[LoadQueue.scala 371:82:@11965.4]
  wire  _T_28346; // @[LoadQueue.scala 371:79:@11966.4]
  wire  _T_28348; // @[LoadQueue.scala 371:82:@11967.4]
  wire  _T_28349; // @[LoadQueue.scala 371:79:@11968.4]
  wire  _T_28351; // @[LoadQueue.scala 371:82:@11969.4]
  wire  _T_28352; // @[LoadQueue.scala 371:79:@11970.4]
  wire  _T_28354; // @[LoadQueue.scala 371:82:@11971.4]
  wire  _T_28355; // @[LoadQueue.scala 371:79:@11972.4]
  wire  _T_28372; // @[LoadQueue.scala 371:96:@11983.4]
  wire  _T_28373; // @[LoadQueue.scala 371:96:@11984.4]
  wire  _T_28374; // @[LoadQueue.scala 371:96:@11985.4]
  wire  _T_28375; // @[LoadQueue.scala 371:96:@11986.4]
  wire  _T_28376; // @[LoadQueue.scala 371:96:@11987.4]
  wire  _T_28377; // @[LoadQueue.scala 371:96:@11988.4]
  assign _GEN_712 = {{2'd0}, tail}; // @[util.scala 14:20:@2870.4]
  assign _T_1020 = 5'h8 - _GEN_712; // @[util.scala 14:20:@2870.4]
  assign _T_1021 = $unsigned(_T_1020); // @[util.scala 14:20:@2871.4]
  assign _T_1022 = _T_1021[4:0]; // @[util.scala 14:20:@2872.4]
  assign _GEN_0 = _T_1022 % 5'h8; // @[util.scala 14:25:@2873.4]
  assign _T_1023 = _GEN_0[3:0]; // @[util.scala 14:25:@2873.4]
  assign _GEN_713 = {{2'd0}, io_bbNumLoads}; // @[LoadQueue.scala 71:46:@2874.4]
  assign _T_1024 = _T_1023 < _GEN_713; // @[LoadQueue.scala 71:46:@2874.4]
  assign initBits_0 = _T_1024 & io_bbStart; // @[LoadQueue.scala 71:63:@2875.4]
  assign _T_1029 = 5'h9 - _GEN_712; // @[util.scala 14:20:@2877.4]
  assign _T_1030 = $unsigned(_T_1029); // @[util.scala 14:20:@2878.4]
  assign _T_1031 = _T_1030[4:0]; // @[util.scala 14:20:@2879.4]
  assign _GEN_8 = _T_1031 % 5'h8; // @[util.scala 14:25:@2880.4]
  assign _T_1032 = _GEN_8[3:0]; // @[util.scala 14:25:@2880.4]
  assign _T_1033 = _T_1032 < _GEN_713; // @[LoadQueue.scala 71:46:@2881.4]
  assign initBits_1 = _T_1033 & io_bbStart; // @[LoadQueue.scala 71:63:@2882.4]
  assign _T_1038 = 5'ha - _GEN_712; // @[util.scala 14:20:@2884.4]
  assign _T_1039 = $unsigned(_T_1038); // @[util.scala 14:20:@2885.4]
  assign _T_1040 = _T_1039[4:0]; // @[util.scala 14:20:@2886.4]
  assign _GEN_18 = _T_1040 % 5'h8; // @[util.scala 14:25:@2887.4]
  assign _T_1041 = _GEN_18[3:0]; // @[util.scala 14:25:@2887.4]
  assign _T_1042 = _T_1041 < _GEN_713; // @[LoadQueue.scala 71:46:@2888.4]
  assign initBits_2 = _T_1042 & io_bbStart; // @[LoadQueue.scala 71:63:@2889.4]
  assign _T_1047 = 5'hb - _GEN_712; // @[util.scala 14:20:@2891.4]
  assign _T_1048 = $unsigned(_T_1047); // @[util.scala 14:20:@2892.4]
  assign _T_1049 = _T_1048[4:0]; // @[util.scala 14:20:@2893.4]
  assign _GEN_26 = _T_1049 % 5'h8; // @[util.scala 14:25:@2894.4]
  assign _T_1050 = _GEN_26[3:0]; // @[util.scala 14:25:@2894.4]
  assign _T_1051 = _T_1050 < _GEN_713; // @[LoadQueue.scala 71:46:@2895.4]
  assign initBits_3 = _T_1051 & io_bbStart; // @[LoadQueue.scala 71:63:@2896.4]
  assign _T_1056 = 5'hc - _GEN_712; // @[util.scala 14:20:@2898.4]
  assign _T_1057 = $unsigned(_T_1056); // @[util.scala 14:20:@2899.4]
  assign _T_1058 = _T_1057[4:0]; // @[util.scala 14:20:@2900.4]
  assign _GEN_36 = _T_1058 % 5'h8; // @[util.scala 14:25:@2901.4]
  assign _T_1059 = _GEN_36[3:0]; // @[util.scala 14:25:@2901.4]
  assign _T_1060 = _T_1059 < _GEN_713; // @[LoadQueue.scala 71:46:@2902.4]
  assign initBits_4 = _T_1060 & io_bbStart; // @[LoadQueue.scala 71:63:@2903.4]
  assign _T_1065 = 5'hd - _GEN_712; // @[util.scala 14:20:@2905.4]
  assign _T_1066 = $unsigned(_T_1065); // @[util.scala 14:20:@2906.4]
  assign _T_1067 = _T_1066[4:0]; // @[util.scala 14:20:@2907.4]
  assign _GEN_44 = _T_1067 % 5'h8; // @[util.scala 14:25:@2908.4]
  assign _T_1068 = _GEN_44[3:0]; // @[util.scala 14:25:@2908.4]
  assign _T_1069 = _T_1068 < _GEN_713; // @[LoadQueue.scala 71:46:@2909.4]
  assign initBits_5 = _T_1069 & io_bbStart; // @[LoadQueue.scala 71:63:@2910.4]
  assign _T_1074 = 5'he - _GEN_712; // @[util.scala 14:20:@2912.4]
  assign _T_1075 = $unsigned(_T_1074); // @[util.scala 14:20:@2913.4]
  assign _T_1076 = _T_1075[4:0]; // @[util.scala 14:20:@2914.4]
  assign _GEN_54 = _T_1076 % 5'h8; // @[util.scala 14:25:@2915.4]
  assign _T_1077 = _GEN_54[3:0]; // @[util.scala 14:25:@2915.4]
  assign _T_1078 = _T_1077 < _GEN_713; // @[LoadQueue.scala 71:46:@2916.4]
  assign initBits_6 = _T_1078 & io_bbStart; // @[LoadQueue.scala 71:63:@2917.4]
  assign _T_1083 = 5'hf - _GEN_712; // @[util.scala 14:20:@2919.4]
  assign _T_1084 = $unsigned(_T_1083); // @[util.scala 14:20:@2920.4]
  assign _T_1085 = _T_1084[4:0]; // @[util.scala 14:20:@2921.4]
  assign _GEN_62 = _T_1085 % 5'h8; // @[util.scala 14:25:@2922.4]
  assign _T_1086 = _GEN_62[3:0]; // @[util.scala 14:25:@2922.4]
  assign _T_1087 = _T_1086 < _GEN_713; // @[LoadQueue.scala 71:46:@2923.4]
  assign initBits_7 = _T_1087 & io_bbStart; // @[LoadQueue.scala 71:63:@2924.4]
  assign _T_1102 = allocatedEntries_0 | initBits_0; // @[LoadQueue.scala 73:78:@2934.4]
  assign _T_1103 = allocatedEntries_1 | initBits_1; // @[LoadQueue.scala 73:78:@2935.4]
  assign _T_1104 = allocatedEntries_2 | initBits_2; // @[LoadQueue.scala 73:78:@2936.4]
  assign _T_1105 = allocatedEntries_3 | initBits_3; // @[LoadQueue.scala 73:78:@2937.4]
  assign _T_1106 = allocatedEntries_4 | initBits_4; // @[LoadQueue.scala 73:78:@2938.4]
  assign _T_1107 = allocatedEntries_5 | initBits_5; // @[LoadQueue.scala 73:78:@2939.4]
  assign _T_1108 = allocatedEntries_6 | initBits_6; // @[LoadQueue.scala 73:78:@2940.4]
  assign _T_1109 = allocatedEntries_7 | initBits_7; // @[LoadQueue.scala 73:78:@2941.4]
  assign _T_1132 = _T_1023[2:0]; // @[:@2965.6]
  assign _GEN_1 = 3'h1 == _T_1132 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2966.6]
  assign _GEN_2 = 3'h2 == _T_1132 ? io_bbLoadOffsets_2 : _GEN_1; // @[LoadQueue.scala 77:20:@2966.6]
  assign _GEN_3 = 3'h3 == _T_1132 ? io_bbLoadOffsets_3 : _GEN_2; // @[LoadQueue.scala 77:20:@2966.6]
  assign _GEN_4 = 3'h4 == _T_1132 ? io_bbLoadOffsets_4 : _GEN_3; // @[LoadQueue.scala 77:20:@2966.6]
  assign _GEN_5 = 3'h5 == _T_1132 ? io_bbLoadOffsets_5 : _GEN_4; // @[LoadQueue.scala 77:20:@2966.6]
  assign _GEN_6 = 3'h6 == _T_1132 ? io_bbLoadOffsets_6 : _GEN_5; // @[LoadQueue.scala 77:20:@2966.6]
  assign _GEN_7 = 3'h7 == _T_1132 ? io_bbLoadOffsets_7 : _GEN_6; // @[LoadQueue.scala 77:20:@2966.6]
  assign _GEN_9 = 3'h1 == _T_1132 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@2973.6]
  assign _GEN_10 = 3'h2 == _T_1132 ? 1'h0 : _GEN_9; // @[LoadQueue.scala 78:18:@2973.6]
  assign _GEN_11 = 3'h3 == _T_1132 ? 1'h0 : _GEN_10; // @[LoadQueue.scala 78:18:@2973.6]
  assign _GEN_12 = 3'h4 == _T_1132 ? 1'h0 : _GEN_11; // @[LoadQueue.scala 78:18:@2973.6]
  assign _GEN_13 = 3'h5 == _T_1132 ? 1'h0 : _GEN_12; // @[LoadQueue.scala 78:18:@2973.6]
  assign _GEN_14 = 3'h6 == _T_1132 ? 1'h0 : _GEN_13; // @[LoadQueue.scala 78:18:@2973.6]
  assign _GEN_15 = 3'h7 == _T_1132 ? 1'h0 : _GEN_14; // @[LoadQueue.scala 78:18:@2973.6]
  assign _GEN_16 = initBits_0 ? _GEN_7 : offsetQ_0; // @[LoadQueue.scala 76:25:@2959.4]
  assign _GEN_17 = initBits_0 ? _GEN_15 : portQ_0; // @[LoadQueue.scala 76:25:@2959.4]
  assign _T_1150 = _T_1032[2:0]; // @[:@2981.6]
  assign _GEN_19 = 3'h1 == _T_1150 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2982.6]
  assign _GEN_20 = 3'h2 == _T_1150 ? io_bbLoadOffsets_2 : _GEN_19; // @[LoadQueue.scala 77:20:@2982.6]
  assign _GEN_21 = 3'h3 == _T_1150 ? io_bbLoadOffsets_3 : _GEN_20; // @[LoadQueue.scala 77:20:@2982.6]
  assign _GEN_22 = 3'h4 == _T_1150 ? io_bbLoadOffsets_4 : _GEN_21; // @[LoadQueue.scala 77:20:@2982.6]
  assign _GEN_23 = 3'h5 == _T_1150 ? io_bbLoadOffsets_5 : _GEN_22; // @[LoadQueue.scala 77:20:@2982.6]
  assign _GEN_24 = 3'h6 == _T_1150 ? io_bbLoadOffsets_6 : _GEN_23; // @[LoadQueue.scala 77:20:@2982.6]
  assign _GEN_25 = 3'h7 == _T_1150 ? io_bbLoadOffsets_7 : _GEN_24; // @[LoadQueue.scala 77:20:@2982.6]
  assign _GEN_27 = 3'h1 == _T_1150 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@2989.6]
  assign _GEN_28 = 3'h2 == _T_1150 ? 1'h0 : _GEN_27; // @[LoadQueue.scala 78:18:@2989.6]
  assign _GEN_29 = 3'h3 == _T_1150 ? 1'h0 : _GEN_28; // @[LoadQueue.scala 78:18:@2989.6]
  assign _GEN_30 = 3'h4 == _T_1150 ? 1'h0 : _GEN_29; // @[LoadQueue.scala 78:18:@2989.6]
  assign _GEN_31 = 3'h5 == _T_1150 ? 1'h0 : _GEN_30; // @[LoadQueue.scala 78:18:@2989.6]
  assign _GEN_32 = 3'h6 == _T_1150 ? 1'h0 : _GEN_31; // @[LoadQueue.scala 78:18:@2989.6]
  assign _GEN_33 = 3'h7 == _T_1150 ? 1'h0 : _GEN_32; // @[LoadQueue.scala 78:18:@2989.6]
  assign _GEN_34 = initBits_1 ? _GEN_25 : offsetQ_1; // @[LoadQueue.scala 76:25:@2975.4]
  assign _GEN_35 = initBits_1 ? _GEN_33 : portQ_1; // @[LoadQueue.scala 76:25:@2975.4]
  assign _T_1168 = _T_1041[2:0]; // @[:@2997.6]
  assign _GEN_37 = 3'h1 == _T_1168 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@2998.6]
  assign _GEN_38 = 3'h2 == _T_1168 ? io_bbLoadOffsets_2 : _GEN_37; // @[LoadQueue.scala 77:20:@2998.6]
  assign _GEN_39 = 3'h3 == _T_1168 ? io_bbLoadOffsets_3 : _GEN_38; // @[LoadQueue.scala 77:20:@2998.6]
  assign _GEN_40 = 3'h4 == _T_1168 ? io_bbLoadOffsets_4 : _GEN_39; // @[LoadQueue.scala 77:20:@2998.6]
  assign _GEN_41 = 3'h5 == _T_1168 ? io_bbLoadOffsets_5 : _GEN_40; // @[LoadQueue.scala 77:20:@2998.6]
  assign _GEN_42 = 3'h6 == _T_1168 ? io_bbLoadOffsets_6 : _GEN_41; // @[LoadQueue.scala 77:20:@2998.6]
  assign _GEN_43 = 3'h7 == _T_1168 ? io_bbLoadOffsets_7 : _GEN_42; // @[LoadQueue.scala 77:20:@2998.6]
  assign _GEN_45 = 3'h1 == _T_1168 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@3005.6]
  assign _GEN_46 = 3'h2 == _T_1168 ? 1'h0 : _GEN_45; // @[LoadQueue.scala 78:18:@3005.6]
  assign _GEN_47 = 3'h3 == _T_1168 ? 1'h0 : _GEN_46; // @[LoadQueue.scala 78:18:@3005.6]
  assign _GEN_48 = 3'h4 == _T_1168 ? 1'h0 : _GEN_47; // @[LoadQueue.scala 78:18:@3005.6]
  assign _GEN_49 = 3'h5 == _T_1168 ? 1'h0 : _GEN_48; // @[LoadQueue.scala 78:18:@3005.6]
  assign _GEN_50 = 3'h6 == _T_1168 ? 1'h0 : _GEN_49; // @[LoadQueue.scala 78:18:@3005.6]
  assign _GEN_51 = 3'h7 == _T_1168 ? 1'h0 : _GEN_50; // @[LoadQueue.scala 78:18:@3005.6]
  assign _GEN_52 = initBits_2 ? _GEN_43 : offsetQ_2; // @[LoadQueue.scala 76:25:@2991.4]
  assign _GEN_53 = initBits_2 ? _GEN_51 : portQ_2; // @[LoadQueue.scala 76:25:@2991.4]
  assign _T_1186 = _T_1050[2:0]; // @[:@3013.6]
  assign _GEN_55 = 3'h1 == _T_1186 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@3014.6]
  assign _GEN_56 = 3'h2 == _T_1186 ? io_bbLoadOffsets_2 : _GEN_55; // @[LoadQueue.scala 77:20:@3014.6]
  assign _GEN_57 = 3'h3 == _T_1186 ? io_bbLoadOffsets_3 : _GEN_56; // @[LoadQueue.scala 77:20:@3014.6]
  assign _GEN_58 = 3'h4 == _T_1186 ? io_bbLoadOffsets_4 : _GEN_57; // @[LoadQueue.scala 77:20:@3014.6]
  assign _GEN_59 = 3'h5 == _T_1186 ? io_bbLoadOffsets_5 : _GEN_58; // @[LoadQueue.scala 77:20:@3014.6]
  assign _GEN_60 = 3'h6 == _T_1186 ? io_bbLoadOffsets_6 : _GEN_59; // @[LoadQueue.scala 77:20:@3014.6]
  assign _GEN_61 = 3'h7 == _T_1186 ? io_bbLoadOffsets_7 : _GEN_60; // @[LoadQueue.scala 77:20:@3014.6]
  assign _GEN_63 = 3'h1 == _T_1186 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@3021.6]
  assign _GEN_64 = 3'h2 == _T_1186 ? 1'h0 : _GEN_63; // @[LoadQueue.scala 78:18:@3021.6]
  assign _GEN_65 = 3'h3 == _T_1186 ? 1'h0 : _GEN_64; // @[LoadQueue.scala 78:18:@3021.6]
  assign _GEN_66 = 3'h4 == _T_1186 ? 1'h0 : _GEN_65; // @[LoadQueue.scala 78:18:@3021.6]
  assign _GEN_67 = 3'h5 == _T_1186 ? 1'h0 : _GEN_66; // @[LoadQueue.scala 78:18:@3021.6]
  assign _GEN_68 = 3'h6 == _T_1186 ? 1'h0 : _GEN_67; // @[LoadQueue.scala 78:18:@3021.6]
  assign _GEN_69 = 3'h7 == _T_1186 ? 1'h0 : _GEN_68; // @[LoadQueue.scala 78:18:@3021.6]
  assign _GEN_70 = initBits_3 ? _GEN_61 : offsetQ_3; // @[LoadQueue.scala 76:25:@3007.4]
  assign _GEN_71 = initBits_3 ? _GEN_69 : portQ_3; // @[LoadQueue.scala 76:25:@3007.4]
  assign _T_1204 = _T_1059[2:0]; // @[:@3029.6]
  assign _GEN_73 = 3'h1 == _T_1204 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@3030.6]
  assign _GEN_74 = 3'h2 == _T_1204 ? io_bbLoadOffsets_2 : _GEN_73; // @[LoadQueue.scala 77:20:@3030.6]
  assign _GEN_75 = 3'h3 == _T_1204 ? io_bbLoadOffsets_3 : _GEN_74; // @[LoadQueue.scala 77:20:@3030.6]
  assign _GEN_76 = 3'h4 == _T_1204 ? io_bbLoadOffsets_4 : _GEN_75; // @[LoadQueue.scala 77:20:@3030.6]
  assign _GEN_77 = 3'h5 == _T_1204 ? io_bbLoadOffsets_5 : _GEN_76; // @[LoadQueue.scala 77:20:@3030.6]
  assign _GEN_78 = 3'h6 == _T_1204 ? io_bbLoadOffsets_6 : _GEN_77; // @[LoadQueue.scala 77:20:@3030.6]
  assign _GEN_79 = 3'h7 == _T_1204 ? io_bbLoadOffsets_7 : _GEN_78; // @[LoadQueue.scala 77:20:@3030.6]
  assign _GEN_81 = 3'h1 == _T_1204 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@3037.6]
  assign _GEN_82 = 3'h2 == _T_1204 ? 1'h0 : _GEN_81; // @[LoadQueue.scala 78:18:@3037.6]
  assign _GEN_83 = 3'h3 == _T_1204 ? 1'h0 : _GEN_82; // @[LoadQueue.scala 78:18:@3037.6]
  assign _GEN_84 = 3'h4 == _T_1204 ? 1'h0 : _GEN_83; // @[LoadQueue.scala 78:18:@3037.6]
  assign _GEN_85 = 3'h5 == _T_1204 ? 1'h0 : _GEN_84; // @[LoadQueue.scala 78:18:@3037.6]
  assign _GEN_86 = 3'h6 == _T_1204 ? 1'h0 : _GEN_85; // @[LoadQueue.scala 78:18:@3037.6]
  assign _GEN_87 = 3'h7 == _T_1204 ? 1'h0 : _GEN_86; // @[LoadQueue.scala 78:18:@3037.6]
  assign _GEN_88 = initBits_4 ? _GEN_79 : offsetQ_4; // @[LoadQueue.scala 76:25:@3023.4]
  assign _GEN_89 = initBits_4 ? _GEN_87 : portQ_4; // @[LoadQueue.scala 76:25:@3023.4]
  assign _T_1222 = _T_1068[2:0]; // @[:@3045.6]
  assign _GEN_91 = 3'h1 == _T_1222 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@3046.6]
  assign _GEN_92 = 3'h2 == _T_1222 ? io_bbLoadOffsets_2 : _GEN_91; // @[LoadQueue.scala 77:20:@3046.6]
  assign _GEN_93 = 3'h3 == _T_1222 ? io_bbLoadOffsets_3 : _GEN_92; // @[LoadQueue.scala 77:20:@3046.6]
  assign _GEN_94 = 3'h4 == _T_1222 ? io_bbLoadOffsets_4 : _GEN_93; // @[LoadQueue.scala 77:20:@3046.6]
  assign _GEN_95 = 3'h5 == _T_1222 ? io_bbLoadOffsets_5 : _GEN_94; // @[LoadQueue.scala 77:20:@3046.6]
  assign _GEN_96 = 3'h6 == _T_1222 ? io_bbLoadOffsets_6 : _GEN_95; // @[LoadQueue.scala 77:20:@3046.6]
  assign _GEN_97 = 3'h7 == _T_1222 ? io_bbLoadOffsets_7 : _GEN_96; // @[LoadQueue.scala 77:20:@3046.6]
  assign _GEN_99 = 3'h1 == _T_1222 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@3053.6]
  assign _GEN_100 = 3'h2 == _T_1222 ? 1'h0 : _GEN_99; // @[LoadQueue.scala 78:18:@3053.6]
  assign _GEN_101 = 3'h3 == _T_1222 ? 1'h0 : _GEN_100; // @[LoadQueue.scala 78:18:@3053.6]
  assign _GEN_102 = 3'h4 == _T_1222 ? 1'h0 : _GEN_101; // @[LoadQueue.scala 78:18:@3053.6]
  assign _GEN_103 = 3'h5 == _T_1222 ? 1'h0 : _GEN_102; // @[LoadQueue.scala 78:18:@3053.6]
  assign _GEN_104 = 3'h6 == _T_1222 ? 1'h0 : _GEN_103; // @[LoadQueue.scala 78:18:@3053.6]
  assign _GEN_105 = 3'h7 == _T_1222 ? 1'h0 : _GEN_104; // @[LoadQueue.scala 78:18:@3053.6]
  assign _GEN_106 = initBits_5 ? _GEN_97 : offsetQ_5; // @[LoadQueue.scala 76:25:@3039.4]
  assign _GEN_107 = initBits_5 ? _GEN_105 : portQ_5; // @[LoadQueue.scala 76:25:@3039.4]
  assign _T_1240 = _T_1077[2:0]; // @[:@3061.6]
  assign _GEN_109 = 3'h1 == _T_1240 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@3062.6]
  assign _GEN_110 = 3'h2 == _T_1240 ? io_bbLoadOffsets_2 : _GEN_109; // @[LoadQueue.scala 77:20:@3062.6]
  assign _GEN_111 = 3'h3 == _T_1240 ? io_bbLoadOffsets_3 : _GEN_110; // @[LoadQueue.scala 77:20:@3062.6]
  assign _GEN_112 = 3'h4 == _T_1240 ? io_bbLoadOffsets_4 : _GEN_111; // @[LoadQueue.scala 77:20:@3062.6]
  assign _GEN_113 = 3'h5 == _T_1240 ? io_bbLoadOffsets_5 : _GEN_112; // @[LoadQueue.scala 77:20:@3062.6]
  assign _GEN_114 = 3'h6 == _T_1240 ? io_bbLoadOffsets_6 : _GEN_113; // @[LoadQueue.scala 77:20:@3062.6]
  assign _GEN_115 = 3'h7 == _T_1240 ? io_bbLoadOffsets_7 : _GEN_114; // @[LoadQueue.scala 77:20:@3062.6]
  assign _GEN_117 = 3'h1 == _T_1240 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@3069.6]
  assign _GEN_118 = 3'h2 == _T_1240 ? 1'h0 : _GEN_117; // @[LoadQueue.scala 78:18:@3069.6]
  assign _GEN_119 = 3'h3 == _T_1240 ? 1'h0 : _GEN_118; // @[LoadQueue.scala 78:18:@3069.6]
  assign _GEN_120 = 3'h4 == _T_1240 ? 1'h0 : _GEN_119; // @[LoadQueue.scala 78:18:@3069.6]
  assign _GEN_121 = 3'h5 == _T_1240 ? 1'h0 : _GEN_120; // @[LoadQueue.scala 78:18:@3069.6]
  assign _GEN_122 = 3'h6 == _T_1240 ? 1'h0 : _GEN_121; // @[LoadQueue.scala 78:18:@3069.6]
  assign _GEN_123 = 3'h7 == _T_1240 ? 1'h0 : _GEN_122; // @[LoadQueue.scala 78:18:@3069.6]
  assign _GEN_124 = initBits_6 ? _GEN_115 : offsetQ_6; // @[LoadQueue.scala 76:25:@3055.4]
  assign _GEN_125 = initBits_6 ? _GEN_123 : portQ_6; // @[LoadQueue.scala 76:25:@3055.4]
  assign _T_1258 = _T_1086[2:0]; // @[:@3077.6]
  assign _GEN_127 = 3'h1 == _T_1258 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@3078.6]
  assign _GEN_128 = 3'h2 == _T_1258 ? io_bbLoadOffsets_2 : _GEN_127; // @[LoadQueue.scala 77:20:@3078.6]
  assign _GEN_129 = 3'h3 == _T_1258 ? io_bbLoadOffsets_3 : _GEN_128; // @[LoadQueue.scala 77:20:@3078.6]
  assign _GEN_130 = 3'h4 == _T_1258 ? io_bbLoadOffsets_4 : _GEN_129; // @[LoadQueue.scala 77:20:@3078.6]
  assign _GEN_131 = 3'h5 == _T_1258 ? io_bbLoadOffsets_5 : _GEN_130; // @[LoadQueue.scala 77:20:@3078.6]
  assign _GEN_132 = 3'h6 == _T_1258 ? io_bbLoadOffsets_6 : _GEN_131; // @[LoadQueue.scala 77:20:@3078.6]
  assign _GEN_133 = 3'h7 == _T_1258 ? io_bbLoadOffsets_7 : _GEN_132; // @[LoadQueue.scala 77:20:@3078.6]
  assign _GEN_135 = 3'h1 == _T_1258 ? io_bbLoadPorts_1 : 1'h0; // @[LoadQueue.scala 78:18:@3085.6]
  assign _GEN_136 = 3'h2 == _T_1258 ? 1'h0 : _GEN_135; // @[LoadQueue.scala 78:18:@3085.6]
  assign _GEN_137 = 3'h3 == _T_1258 ? 1'h0 : _GEN_136; // @[LoadQueue.scala 78:18:@3085.6]
  assign _GEN_138 = 3'h4 == _T_1258 ? 1'h0 : _GEN_137; // @[LoadQueue.scala 78:18:@3085.6]
  assign _GEN_139 = 3'h5 == _T_1258 ? 1'h0 : _GEN_138; // @[LoadQueue.scala 78:18:@3085.6]
  assign _GEN_140 = 3'h6 == _T_1258 ? 1'h0 : _GEN_139; // @[LoadQueue.scala 78:18:@3085.6]
  assign _GEN_141 = 3'h7 == _T_1258 ? 1'h0 : _GEN_140; // @[LoadQueue.scala 78:18:@3085.6]
  assign _GEN_142 = initBits_7 ? _GEN_133 : offsetQ_7; // @[LoadQueue.scala 76:25:@3071.4]
  assign _GEN_143 = initBits_7 ? _GEN_141 : portQ_7; // @[LoadQueue.scala 76:25:@3071.4]
  assign _T_1280 = _GEN_7 + 3'h1; // @[util.scala 10:8:@3096.6]
  assign _GEN_72 = _T_1280 % 4'h8; // @[util.scala 10:14:@3097.6]
  assign _T_1281 = _GEN_72[3:0]; // @[util.scala 10:14:@3097.6]
  assign _GEN_745 = {{1'd0}, io_storeTail}; // @[LoadQueue.scala 97:56:@3098.6]
  assign _T_1282 = _T_1281 == _GEN_745; // @[LoadQueue.scala 97:56:@3098.6]
  assign _T_1283 = io_storeEmpty & _T_1282; // @[LoadQueue.scala 96:50:@3099.6]
  assign _T_1285 = _T_1283 == 1'h0; // @[LoadQueue.scala 96:34:@3100.6]
  assign _T_1287 = previousStoreHead <= offsetQ_0; // @[LoadQueue.scala 101:36:@3108.8]
  assign _T_1288 = offsetQ_0 < io_storeHead; // @[LoadQueue.scala 101:86:@3109.8]
  assign _T_1289 = _T_1287 & _T_1288; // @[LoadQueue.scala 101:61:@3110.8]
  assign _T_1291 = previousStoreHead > io_storeHead; // @[LoadQueue.scala 103:36:@3115.10]
  assign _T_1292 = io_storeHead <= offsetQ_0; // @[LoadQueue.scala 103:69:@3116.10]
  assign _T_1293 = offsetQ_0 < previousStoreHead; // @[LoadQueue.scala 104:31:@3117.10]
  assign _T_1294 = _T_1292 & _T_1293; // @[LoadQueue.scala 103:94:@3118.10]
  assign _T_1296 = _T_1294 == 1'h0; // @[LoadQueue.scala 103:54:@3119.10]
  assign _T_1297 = _T_1291 & _T_1296; // @[LoadQueue.scala 103:51:@3120.10]
  assign _GEN_152 = _T_1297 ? 1'h0 : checkBits_0; // @[LoadQueue.scala 104:53:@3121.10]
  assign _GEN_153 = _T_1289 ? 1'h0 : _GEN_152; // @[LoadQueue.scala 101:102:@3111.8]
  assign _GEN_154 = io_storeEmpty ? 1'h0 : _GEN_153; // @[LoadQueue.scala 99:27:@3104.6]
  assign _GEN_155 = initBits_0 ? _T_1285 : _GEN_154; // @[LoadQueue.scala 95:34:@3089.4]
  assign _T_1310 = _GEN_25 + 3'h1; // @[util.scala 10:8:@3132.6]
  assign _GEN_80 = _T_1310 % 4'h8; // @[util.scala 10:14:@3133.6]
  assign _T_1311 = _GEN_80[3:0]; // @[util.scala 10:14:@3133.6]
  assign _T_1312 = _T_1311 == _GEN_745; // @[LoadQueue.scala 97:56:@3134.6]
  assign _T_1313 = io_storeEmpty & _T_1312; // @[LoadQueue.scala 96:50:@3135.6]
  assign _T_1315 = _T_1313 == 1'h0; // @[LoadQueue.scala 96:34:@3136.6]
  assign _T_1317 = previousStoreHead <= offsetQ_1; // @[LoadQueue.scala 101:36:@3144.8]
  assign _T_1318 = offsetQ_1 < io_storeHead; // @[LoadQueue.scala 101:86:@3145.8]
  assign _T_1319 = _T_1317 & _T_1318; // @[LoadQueue.scala 101:61:@3146.8]
  assign _T_1322 = io_storeHead <= offsetQ_1; // @[LoadQueue.scala 103:69:@3152.10]
  assign _T_1323 = offsetQ_1 < previousStoreHead; // @[LoadQueue.scala 104:31:@3153.10]
  assign _T_1324 = _T_1322 & _T_1323; // @[LoadQueue.scala 103:94:@3154.10]
  assign _T_1326 = _T_1324 == 1'h0; // @[LoadQueue.scala 103:54:@3155.10]
  assign _T_1327 = _T_1291 & _T_1326; // @[LoadQueue.scala 103:51:@3156.10]
  assign _GEN_164 = _T_1327 ? 1'h0 : checkBits_1; // @[LoadQueue.scala 104:53:@3157.10]
  assign _GEN_165 = _T_1319 ? 1'h0 : _GEN_164; // @[LoadQueue.scala 101:102:@3147.8]
  assign _GEN_166 = io_storeEmpty ? 1'h0 : _GEN_165; // @[LoadQueue.scala 99:27:@3140.6]
  assign _GEN_167 = initBits_1 ? _T_1315 : _GEN_166; // @[LoadQueue.scala 95:34:@3125.4]
  assign _T_1340 = _GEN_43 + 3'h1; // @[util.scala 10:8:@3168.6]
  assign _GEN_90 = _T_1340 % 4'h8; // @[util.scala 10:14:@3169.6]
  assign _T_1341 = _GEN_90[3:0]; // @[util.scala 10:14:@3169.6]
  assign _T_1342 = _T_1341 == _GEN_745; // @[LoadQueue.scala 97:56:@3170.6]
  assign _T_1343 = io_storeEmpty & _T_1342; // @[LoadQueue.scala 96:50:@3171.6]
  assign _T_1345 = _T_1343 == 1'h0; // @[LoadQueue.scala 96:34:@3172.6]
  assign _T_1347 = previousStoreHead <= offsetQ_2; // @[LoadQueue.scala 101:36:@3180.8]
  assign _T_1348 = offsetQ_2 < io_storeHead; // @[LoadQueue.scala 101:86:@3181.8]
  assign _T_1349 = _T_1347 & _T_1348; // @[LoadQueue.scala 101:61:@3182.8]
  assign _T_1352 = io_storeHead <= offsetQ_2; // @[LoadQueue.scala 103:69:@3188.10]
  assign _T_1353 = offsetQ_2 < previousStoreHead; // @[LoadQueue.scala 104:31:@3189.10]
  assign _T_1354 = _T_1352 & _T_1353; // @[LoadQueue.scala 103:94:@3190.10]
  assign _T_1356 = _T_1354 == 1'h0; // @[LoadQueue.scala 103:54:@3191.10]
  assign _T_1357 = _T_1291 & _T_1356; // @[LoadQueue.scala 103:51:@3192.10]
  assign _GEN_176 = _T_1357 ? 1'h0 : checkBits_2; // @[LoadQueue.scala 104:53:@3193.10]
  assign _GEN_177 = _T_1349 ? 1'h0 : _GEN_176; // @[LoadQueue.scala 101:102:@3183.8]
  assign _GEN_178 = io_storeEmpty ? 1'h0 : _GEN_177; // @[LoadQueue.scala 99:27:@3176.6]
  assign _GEN_179 = initBits_2 ? _T_1345 : _GEN_178; // @[LoadQueue.scala 95:34:@3161.4]
  assign _T_1370 = _GEN_61 + 3'h1; // @[util.scala 10:8:@3204.6]
  assign _GEN_98 = _T_1370 % 4'h8; // @[util.scala 10:14:@3205.6]
  assign _T_1371 = _GEN_98[3:0]; // @[util.scala 10:14:@3205.6]
  assign _T_1372 = _T_1371 == _GEN_745; // @[LoadQueue.scala 97:56:@3206.6]
  assign _T_1373 = io_storeEmpty & _T_1372; // @[LoadQueue.scala 96:50:@3207.6]
  assign _T_1375 = _T_1373 == 1'h0; // @[LoadQueue.scala 96:34:@3208.6]
  assign _T_1377 = previousStoreHead <= offsetQ_3; // @[LoadQueue.scala 101:36:@3216.8]
  assign _T_1378 = offsetQ_3 < io_storeHead; // @[LoadQueue.scala 101:86:@3217.8]
  assign _T_1379 = _T_1377 & _T_1378; // @[LoadQueue.scala 101:61:@3218.8]
  assign _T_1382 = io_storeHead <= offsetQ_3; // @[LoadQueue.scala 103:69:@3224.10]
  assign _T_1383 = offsetQ_3 < previousStoreHead; // @[LoadQueue.scala 104:31:@3225.10]
  assign _T_1384 = _T_1382 & _T_1383; // @[LoadQueue.scala 103:94:@3226.10]
  assign _T_1386 = _T_1384 == 1'h0; // @[LoadQueue.scala 103:54:@3227.10]
  assign _T_1387 = _T_1291 & _T_1386; // @[LoadQueue.scala 103:51:@3228.10]
  assign _GEN_188 = _T_1387 ? 1'h0 : checkBits_3; // @[LoadQueue.scala 104:53:@3229.10]
  assign _GEN_189 = _T_1379 ? 1'h0 : _GEN_188; // @[LoadQueue.scala 101:102:@3219.8]
  assign _GEN_190 = io_storeEmpty ? 1'h0 : _GEN_189; // @[LoadQueue.scala 99:27:@3212.6]
  assign _GEN_191 = initBits_3 ? _T_1375 : _GEN_190; // @[LoadQueue.scala 95:34:@3197.4]
  assign _T_1400 = _GEN_79 + 3'h1; // @[util.scala 10:8:@3240.6]
  assign _GEN_108 = _T_1400 % 4'h8; // @[util.scala 10:14:@3241.6]
  assign _T_1401 = _GEN_108[3:0]; // @[util.scala 10:14:@3241.6]
  assign _T_1402 = _T_1401 == _GEN_745; // @[LoadQueue.scala 97:56:@3242.6]
  assign _T_1403 = io_storeEmpty & _T_1402; // @[LoadQueue.scala 96:50:@3243.6]
  assign _T_1405 = _T_1403 == 1'h0; // @[LoadQueue.scala 96:34:@3244.6]
  assign _T_1407 = previousStoreHead <= offsetQ_4; // @[LoadQueue.scala 101:36:@3252.8]
  assign _T_1408 = offsetQ_4 < io_storeHead; // @[LoadQueue.scala 101:86:@3253.8]
  assign _T_1409 = _T_1407 & _T_1408; // @[LoadQueue.scala 101:61:@3254.8]
  assign _T_1412 = io_storeHead <= offsetQ_4; // @[LoadQueue.scala 103:69:@3260.10]
  assign _T_1413 = offsetQ_4 < previousStoreHead; // @[LoadQueue.scala 104:31:@3261.10]
  assign _T_1414 = _T_1412 & _T_1413; // @[LoadQueue.scala 103:94:@3262.10]
  assign _T_1416 = _T_1414 == 1'h0; // @[LoadQueue.scala 103:54:@3263.10]
  assign _T_1417 = _T_1291 & _T_1416; // @[LoadQueue.scala 103:51:@3264.10]
  assign _GEN_200 = _T_1417 ? 1'h0 : checkBits_4; // @[LoadQueue.scala 104:53:@3265.10]
  assign _GEN_201 = _T_1409 ? 1'h0 : _GEN_200; // @[LoadQueue.scala 101:102:@3255.8]
  assign _GEN_202 = io_storeEmpty ? 1'h0 : _GEN_201; // @[LoadQueue.scala 99:27:@3248.6]
  assign _GEN_203 = initBits_4 ? _T_1405 : _GEN_202; // @[LoadQueue.scala 95:34:@3233.4]
  assign _T_1430 = _GEN_97 + 3'h1; // @[util.scala 10:8:@3276.6]
  assign _GEN_116 = _T_1430 % 4'h8; // @[util.scala 10:14:@3277.6]
  assign _T_1431 = _GEN_116[3:0]; // @[util.scala 10:14:@3277.6]
  assign _T_1432 = _T_1431 == _GEN_745; // @[LoadQueue.scala 97:56:@3278.6]
  assign _T_1433 = io_storeEmpty & _T_1432; // @[LoadQueue.scala 96:50:@3279.6]
  assign _T_1435 = _T_1433 == 1'h0; // @[LoadQueue.scala 96:34:@3280.6]
  assign _T_1437 = previousStoreHead <= offsetQ_5; // @[LoadQueue.scala 101:36:@3288.8]
  assign _T_1438 = offsetQ_5 < io_storeHead; // @[LoadQueue.scala 101:86:@3289.8]
  assign _T_1439 = _T_1437 & _T_1438; // @[LoadQueue.scala 101:61:@3290.8]
  assign _T_1442 = io_storeHead <= offsetQ_5; // @[LoadQueue.scala 103:69:@3296.10]
  assign _T_1443 = offsetQ_5 < previousStoreHead; // @[LoadQueue.scala 104:31:@3297.10]
  assign _T_1444 = _T_1442 & _T_1443; // @[LoadQueue.scala 103:94:@3298.10]
  assign _T_1446 = _T_1444 == 1'h0; // @[LoadQueue.scala 103:54:@3299.10]
  assign _T_1447 = _T_1291 & _T_1446; // @[LoadQueue.scala 103:51:@3300.10]
  assign _GEN_212 = _T_1447 ? 1'h0 : checkBits_5; // @[LoadQueue.scala 104:53:@3301.10]
  assign _GEN_213 = _T_1439 ? 1'h0 : _GEN_212; // @[LoadQueue.scala 101:102:@3291.8]
  assign _GEN_214 = io_storeEmpty ? 1'h0 : _GEN_213; // @[LoadQueue.scala 99:27:@3284.6]
  assign _GEN_215 = initBits_5 ? _T_1435 : _GEN_214; // @[LoadQueue.scala 95:34:@3269.4]
  assign _T_1460 = _GEN_115 + 3'h1; // @[util.scala 10:8:@3312.6]
  assign _GEN_126 = _T_1460 % 4'h8; // @[util.scala 10:14:@3313.6]
  assign _T_1461 = _GEN_126[3:0]; // @[util.scala 10:14:@3313.6]
  assign _T_1462 = _T_1461 == _GEN_745; // @[LoadQueue.scala 97:56:@3314.6]
  assign _T_1463 = io_storeEmpty & _T_1462; // @[LoadQueue.scala 96:50:@3315.6]
  assign _T_1465 = _T_1463 == 1'h0; // @[LoadQueue.scala 96:34:@3316.6]
  assign _T_1467 = previousStoreHead <= offsetQ_6; // @[LoadQueue.scala 101:36:@3324.8]
  assign _T_1468 = offsetQ_6 < io_storeHead; // @[LoadQueue.scala 101:86:@3325.8]
  assign _T_1469 = _T_1467 & _T_1468; // @[LoadQueue.scala 101:61:@3326.8]
  assign _T_1472 = io_storeHead <= offsetQ_6; // @[LoadQueue.scala 103:69:@3332.10]
  assign _T_1473 = offsetQ_6 < previousStoreHead; // @[LoadQueue.scala 104:31:@3333.10]
  assign _T_1474 = _T_1472 & _T_1473; // @[LoadQueue.scala 103:94:@3334.10]
  assign _T_1476 = _T_1474 == 1'h0; // @[LoadQueue.scala 103:54:@3335.10]
  assign _T_1477 = _T_1291 & _T_1476; // @[LoadQueue.scala 103:51:@3336.10]
  assign _GEN_224 = _T_1477 ? 1'h0 : checkBits_6; // @[LoadQueue.scala 104:53:@3337.10]
  assign _GEN_225 = _T_1469 ? 1'h0 : _GEN_224; // @[LoadQueue.scala 101:102:@3327.8]
  assign _GEN_226 = io_storeEmpty ? 1'h0 : _GEN_225; // @[LoadQueue.scala 99:27:@3320.6]
  assign _GEN_227 = initBits_6 ? _T_1465 : _GEN_226; // @[LoadQueue.scala 95:34:@3305.4]
  assign _T_1490 = _GEN_133 + 3'h1; // @[util.scala 10:8:@3348.6]
  assign _GEN_134 = _T_1490 % 4'h8; // @[util.scala 10:14:@3349.6]
  assign _T_1491 = _GEN_134[3:0]; // @[util.scala 10:14:@3349.6]
  assign _T_1492 = _T_1491 == _GEN_745; // @[LoadQueue.scala 97:56:@3350.6]
  assign _T_1493 = io_storeEmpty & _T_1492; // @[LoadQueue.scala 96:50:@3351.6]
  assign _T_1495 = _T_1493 == 1'h0; // @[LoadQueue.scala 96:34:@3352.6]
  assign _T_1497 = previousStoreHead <= offsetQ_7; // @[LoadQueue.scala 101:36:@3360.8]
  assign _T_1498 = offsetQ_7 < io_storeHead; // @[LoadQueue.scala 101:86:@3361.8]
  assign _T_1499 = _T_1497 & _T_1498; // @[LoadQueue.scala 101:61:@3362.8]
  assign _T_1502 = io_storeHead <= offsetQ_7; // @[LoadQueue.scala 103:69:@3368.10]
  assign _T_1503 = offsetQ_7 < previousStoreHead; // @[LoadQueue.scala 104:31:@3369.10]
  assign _T_1504 = _T_1502 & _T_1503; // @[LoadQueue.scala 103:94:@3370.10]
  assign _T_1506 = _T_1504 == 1'h0; // @[LoadQueue.scala 103:54:@3371.10]
  assign _T_1507 = _T_1291 & _T_1506; // @[LoadQueue.scala 103:51:@3372.10]
  assign _GEN_236 = _T_1507 ? 1'h0 : checkBits_7; // @[LoadQueue.scala 104:53:@3373.10]
  assign _GEN_237 = _T_1499 ? 1'h0 : _GEN_236; // @[LoadQueue.scala 101:102:@3363.8]
  assign _GEN_238 = io_storeEmpty ? 1'h0 : _GEN_237; // @[LoadQueue.scala 99:27:@3356.6]
  assign _GEN_239 = initBits_7 ? _T_1495 : _GEN_238; // @[LoadQueue.scala 95:34:@3341.4]
  assign _T_1511 = 8'h1 << io_storeHead; // @[OneHot.scala 52:12:@3378.4]
  assign _T_1513 = _T_1511[0]; // @[util.scala 60:60:@3380.4]
  assign _T_1514 = _T_1511[1]; // @[util.scala 60:60:@3381.4]
  assign _T_1515 = _T_1511[2]; // @[util.scala 60:60:@3382.4]
  assign _T_1516 = _T_1511[3]; // @[util.scala 60:60:@3383.4]
  assign _T_1517 = _T_1511[4]; // @[util.scala 60:60:@3384.4]
  assign _T_1518 = _T_1511[5]; // @[util.scala 60:60:@3385.4]
  assign _T_1519 = _T_1511[6]; // @[util.scala 60:60:@3386.4]
  assign _T_1520 = _T_1511[7]; // @[util.scala 60:60:@3387.4]
  assign _T_2299 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0}; // @[Mux.scala 19:72:@3839.4]
  assign _T_2301 = _T_1513 ? _T_2299 : 256'h0; // @[Mux.scala 19:72:@3840.4]
  assign _T_2308 = {io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1}; // @[Mux.scala 19:72:@3847.4]
  assign _T_2310 = _T_1514 ? _T_2308 : 256'h0; // @[Mux.scala 19:72:@3848.4]
  assign _T_2317 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2}; // @[Mux.scala 19:72:@3855.4]
  assign _T_2319 = _T_1515 ? _T_2317 : 256'h0; // @[Mux.scala 19:72:@3856.4]
  assign _T_2326 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3}; // @[Mux.scala 19:72:@3863.4]
  assign _T_2328 = _T_1516 ? _T_2326 : 256'h0; // @[Mux.scala 19:72:@3864.4]
  assign _T_2335 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4}; // @[Mux.scala 19:72:@3871.4]
  assign _T_2337 = _T_1517 ? _T_2335 : 256'h0; // @[Mux.scala 19:72:@3872.4]
  assign _T_2344 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5}; // @[Mux.scala 19:72:@3879.4]
  assign _T_2346 = _T_1518 ? _T_2344 : 256'h0; // @[Mux.scala 19:72:@3880.4]
  assign _T_2353 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7,io_storeDataQueue_6}; // @[Mux.scala 19:72:@3887.4]
  assign _T_2355 = _T_1519 ? _T_2353 : 256'h0; // @[Mux.scala 19:72:@3888.4]
  assign _T_2362 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_7}; // @[Mux.scala 19:72:@3895.4]
  assign _T_2364 = _T_1520 ? _T_2362 : 256'h0; // @[Mux.scala 19:72:@3896.4]
  assign _T_2365 = _T_2301 | _T_2310; // @[Mux.scala 19:72:@3897.4]
  assign _T_2366 = _T_2365 | _T_2319; // @[Mux.scala 19:72:@3898.4]
  assign _T_2367 = _T_2366 | _T_2328; // @[Mux.scala 19:72:@3899.4]
  assign _T_2368 = _T_2367 | _T_2337; // @[Mux.scala 19:72:@3900.4]
  assign _T_2369 = _T_2368 | _T_2346; // @[Mux.scala 19:72:@3901.4]
  assign _T_2370 = _T_2369 | _T_2355; // @[Mux.scala 19:72:@3902.4]
  assign _T_2371 = _T_2370 | _T_2364; // @[Mux.scala 19:72:@3903.4]
  assign _T_2612 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0}; // @[Mux.scala 19:72:@4021.4]
  assign _T_2614 = _T_1513 ? _T_2612 : 8'h0; // @[Mux.scala 19:72:@4022.4]
  assign _T_2621 = {io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1}; // @[Mux.scala 19:72:@4029.4]
  assign _T_2623 = _T_1514 ? _T_2621 : 8'h0; // @[Mux.scala 19:72:@4030.4]
  assign _T_2630 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2}; // @[Mux.scala 19:72:@4037.4]
  assign _T_2632 = _T_1515 ? _T_2630 : 8'h0; // @[Mux.scala 19:72:@4038.4]
  assign _T_2639 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3}; // @[Mux.scala 19:72:@4045.4]
  assign _T_2641 = _T_1516 ? _T_2639 : 8'h0; // @[Mux.scala 19:72:@4046.4]
  assign _T_2648 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4}; // @[Mux.scala 19:72:@4053.4]
  assign _T_2650 = _T_1517 ? _T_2648 : 8'h0; // @[Mux.scala 19:72:@4054.4]
  assign _T_2657 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5}; // @[Mux.scala 19:72:@4061.4]
  assign _T_2659 = _T_1518 ? _T_2657 : 8'h0; // @[Mux.scala 19:72:@4062.4]
  assign _T_2666 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7,io_storeDataDone_6}; // @[Mux.scala 19:72:@4069.4]
  assign _T_2668 = _T_1519 ? _T_2666 : 8'h0; // @[Mux.scala 19:72:@4070.4]
  assign _T_2675 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_7}; // @[Mux.scala 19:72:@4077.4]
  assign _T_2677 = _T_1520 ? _T_2675 : 8'h0; // @[Mux.scala 19:72:@4078.4]
  assign _T_2678 = _T_2614 | _T_2623; // @[Mux.scala 19:72:@4079.4]
  assign _T_2679 = _T_2678 | _T_2632; // @[Mux.scala 19:72:@4080.4]
  assign _T_2680 = _T_2679 | _T_2641; // @[Mux.scala 19:72:@4081.4]
  assign _T_2681 = _T_2680 | _T_2650; // @[Mux.scala 19:72:@4082.4]
  assign _T_2682 = _T_2681 | _T_2659; // @[Mux.scala 19:72:@4083.4]
  assign _T_2683 = _T_2682 | _T_2668; // @[Mux.scala 19:72:@4084.4]
  assign _T_2684 = _T_2683 | _T_2677; // @[Mux.scala 19:72:@4085.4]
  assign _T_2761 = io_storeHead < io_storeTail; // @[LoadQueue.scala 121:105:@4105.4]
  assign _T_2763 = io_storeHead <= 3'h0; // @[LoadQueue.scala 122:18:@4106.4]
  assign _T_2765 = 3'h0 < io_storeTail; // @[LoadQueue.scala 122:36:@4107.4]
  assign _T_2766 = _T_2763 & _T_2765; // @[LoadQueue.scala 122:27:@4108.4]
  assign _T_2768 = io_storeEmpty == 1'h0; // @[LoadQueue.scala 122:52:@4109.4]
  assign _T_2770 = io_storeTail <= 3'h0; // @[LoadQueue.scala 122:85:@4110.4]
  assign _T_2772 = 3'h0 < io_storeHead; // @[LoadQueue.scala 122:103:@4111.4]
  assign _T_2773 = _T_2770 & _T_2772; // @[LoadQueue.scala 122:94:@4112.4]
  assign _T_2775 = _T_2773 == 1'h0; // @[LoadQueue.scala 122:70:@4113.4]
  assign _T_2776 = _T_2768 & _T_2775; // @[LoadQueue.scala 122:67:@4114.4]
  assign validEntriesInStoreQ_0 = _T_2761 ? _T_2766 : _T_2776; // @[LoadQueue.scala 121:91:@4115.4]
  assign _T_2780 = io_storeHead <= 3'h1; // @[LoadQueue.scala 122:18:@4117.4]
  assign _T_2782 = 3'h1 < io_storeTail; // @[LoadQueue.scala 122:36:@4118.4]
  assign _T_2783 = _T_2780 & _T_2782; // @[LoadQueue.scala 122:27:@4119.4]
  assign _T_2787 = io_storeTail <= 3'h1; // @[LoadQueue.scala 122:85:@4121.4]
  assign _T_2789 = 3'h1 < io_storeHead; // @[LoadQueue.scala 122:103:@4122.4]
  assign _T_2790 = _T_2787 & _T_2789; // @[LoadQueue.scala 122:94:@4123.4]
  assign _T_2792 = _T_2790 == 1'h0; // @[LoadQueue.scala 122:70:@4124.4]
  assign _T_2793 = _T_2768 & _T_2792; // @[LoadQueue.scala 122:67:@4125.4]
  assign validEntriesInStoreQ_1 = _T_2761 ? _T_2783 : _T_2793; // @[LoadQueue.scala 121:91:@4126.4]
  assign _T_2797 = io_storeHead <= 3'h2; // @[LoadQueue.scala 122:18:@4128.4]
  assign _T_2799 = 3'h2 < io_storeTail; // @[LoadQueue.scala 122:36:@4129.4]
  assign _T_2800 = _T_2797 & _T_2799; // @[LoadQueue.scala 122:27:@4130.4]
  assign _T_2804 = io_storeTail <= 3'h2; // @[LoadQueue.scala 122:85:@4132.4]
  assign _T_2806 = 3'h2 < io_storeHead; // @[LoadQueue.scala 122:103:@4133.4]
  assign _T_2807 = _T_2804 & _T_2806; // @[LoadQueue.scala 122:94:@4134.4]
  assign _T_2809 = _T_2807 == 1'h0; // @[LoadQueue.scala 122:70:@4135.4]
  assign _T_2810 = _T_2768 & _T_2809; // @[LoadQueue.scala 122:67:@4136.4]
  assign validEntriesInStoreQ_2 = _T_2761 ? _T_2800 : _T_2810; // @[LoadQueue.scala 121:91:@4137.4]
  assign _T_2814 = io_storeHead <= 3'h3; // @[LoadQueue.scala 122:18:@4139.4]
  assign _T_2816 = 3'h3 < io_storeTail; // @[LoadQueue.scala 122:36:@4140.4]
  assign _T_2817 = _T_2814 & _T_2816; // @[LoadQueue.scala 122:27:@4141.4]
  assign _T_2821 = io_storeTail <= 3'h3; // @[LoadQueue.scala 122:85:@4143.4]
  assign _T_2823 = 3'h3 < io_storeHead; // @[LoadQueue.scala 122:103:@4144.4]
  assign _T_2824 = _T_2821 & _T_2823; // @[LoadQueue.scala 122:94:@4145.4]
  assign _T_2826 = _T_2824 == 1'h0; // @[LoadQueue.scala 122:70:@4146.4]
  assign _T_2827 = _T_2768 & _T_2826; // @[LoadQueue.scala 122:67:@4147.4]
  assign validEntriesInStoreQ_3 = _T_2761 ? _T_2817 : _T_2827; // @[LoadQueue.scala 121:91:@4148.4]
  assign _T_2831 = io_storeHead <= 3'h4; // @[LoadQueue.scala 122:18:@4150.4]
  assign _T_2833 = 3'h4 < io_storeTail; // @[LoadQueue.scala 122:36:@4151.4]
  assign _T_2834 = _T_2831 & _T_2833; // @[LoadQueue.scala 122:27:@4152.4]
  assign _T_2838 = io_storeTail <= 3'h4; // @[LoadQueue.scala 122:85:@4154.4]
  assign _T_2840 = 3'h4 < io_storeHead; // @[LoadQueue.scala 122:103:@4155.4]
  assign _T_2841 = _T_2838 & _T_2840; // @[LoadQueue.scala 122:94:@4156.4]
  assign _T_2843 = _T_2841 == 1'h0; // @[LoadQueue.scala 122:70:@4157.4]
  assign _T_2844 = _T_2768 & _T_2843; // @[LoadQueue.scala 122:67:@4158.4]
  assign validEntriesInStoreQ_4 = _T_2761 ? _T_2834 : _T_2844; // @[LoadQueue.scala 121:91:@4159.4]
  assign _T_2848 = io_storeHead <= 3'h5; // @[LoadQueue.scala 122:18:@4161.4]
  assign _T_2850 = 3'h5 < io_storeTail; // @[LoadQueue.scala 122:36:@4162.4]
  assign _T_2851 = _T_2848 & _T_2850; // @[LoadQueue.scala 122:27:@4163.4]
  assign _T_2855 = io_storeTail <= 3'h5; // @[LoadQueue.scala 122:85:@4165.4]
  assign _T_2857 = 3'h5 < io_storeHead; // @[LoadQueue.scala 122:103:@4166.4]
  assign _T_2858 = _T_2855 & _T_2857; // @[LoadQueue.scala 122:94:@4167.4]
  assign _T_2860 = _T_2858 == 1'h0; // @[LoadQueue.scala 122:70:@4168.4]
  assign _T_2861 = _T_2768 & _T_2860; // @[LoadQueue.scala 122:67:@4169.4]
  assign validEntriesInStoreQ_5 = _T_2761 ? _T_2851 : _T_2861; // @[LoadQueue.scala 121:91:@4170.4]
  assign _T_2865 = io_storeHead <= 3'h6; // @[LoadQueue.scala 122:18:@4172.4]
  assign _T_2867 = 3'h6 < io_storeTail; // @[LoadQueue.scala 122:36:@4173.4]
  assign _T_2868 = _T_2865 & _T_2867; // @[LoadQueue.scala 122:27:@4174.4]
  assign _T_2872 = io_storeTail <= 3'h6; // @[LoadQueue.scala 122:85:@4176.4]
  assign _T_2874 = 3'h6 < io_storeHead; // @[LoadQueue.scala 122:103:@4177.4]
  assign _T_2875 = _T_2872 & _T_2874; // @[LoadQueue.scala 122:94:@4178.4]
  assign _T_2877 = _T_2875 == 1'h0; // @[LoadQueue.scala 122:70:@4179.4]
  assign _T_2878 = _T_2768 & _T_2877; // @[LoadQueue.scala 122:67:@4180.4]
  assign validEntriesInStoreQ_6 = _T_2761 ? _T_2868 : _T_2878; // @[LoadQueue.scala 121:91:@4181.4]
  assign validEntriesInStoreQ_7 = _T_2761 ? 1'h0 : _T_2768; // @[LoadQueue.scala 121:91:@4192.4]
  assign storesToCheck_0_0 = _T_1292 ? _T_2763 : 1'h1; // @[LoadQueue.scala 131:10:@4211.4]
  assign _T_3294 = 3'h1 <= offsetQ_0; // @[LoadQueue.scala 131:81:@4214.4]
  assign _T_3295 = _T_2780 & _T_3294; // @[LoadQueue.scala 131:72:@4215.4]
  assign _T_3297 = offsetQ_0 < 3'h1; // @[LoadQueue.scala 132:33:@4216.4]
  assign _T_3300 = _T_3297 & _T_2789; // @[LoadQueue.scala 132:41:@4218.4]
  assign _T_3302 = _T_3300 == 1'h0; // @[LoadQueue.scala 132:9:@4219.4]
  assign storesToCheck_0_1 = _T_1292 ? _T_3295 : _T_3302; // @[LoadQueue.scala 131:10:@4220.4]
  assign _T_3308 = 3'h2 <= offsetQ_0; // @[LoadQueue.scala 131:81:@4223.4]
  assign _T_3309 = _T_2797 & _T_3308; // @[LoadQueue.scala 131:72:@4224.4]
  assign _T_3311 = offsetQ_0 < 3'h2; // @[LoadQueue.scala 132:33:@4225.4]
  assign _T_3314 = _T_3311 & _T_2806; // @[LoadQueue.scala 132:41:@4227.4]
  assign _T_3316 = _T_3314 == 1'h0; // @[LoadQueue.scala 132:9:@4228.4]
  assign storesToCheck_0_2 = _T_1292 ? _T_3309 : _T_3316; // @[LoadQueue.scala 131:10:@4229.4]
  assign _T_3322 = 3'h3 <= offsetQ_0; // @[LoadQueue.scala 131:81:@4232.4]
  assign _T_3323 = _T_2814 & _T_3322; // @[LoadQueue.scala 131:72:@4233.4]
  assign _T_3325 = offsetQ_0 < 3'h3; // @[LoadQueue.scala 132:33:@4234.4]
  assign _T_3328 = _T_3325 & _T_2823; // @[LoadQueue.scala 132:41:@4236.4]
  assign _T_3330 = _T_3328 == 1'h0; // @[LoadQueue.scala 132:9:@4237.4]
  assign storesToCheck_0_3 = _T_1292 ? _T_3323 : _T_3330; // @[LoadQueue.scala 131:10:@4238.4]
  assign _T_3336 = 3'h4 <= offsetQ_0; // @[LoadQueue.scala 131:81:@4241.4]
  assign _T_3337 = _T_2831 & _T_3336; // @[LoadQueue.scala 131:72:@4242.4]
  assign _T_3339 = offsetQ_0 < 3'h4; // @[LoadQueue.scala 132:33:@4243.4]
  assign _T_3342 = _T_3339 & _T_2840; // @[LoadQueue.scala 132:41:@4245.4]
  assign _T_3344 = _T_3342 == 1'h0; // @[LoadQueue.scala 132:9:@4246.4]
  assign storesToCheck_0_4 = _T_1292 ? _T_3337 : _T_3344; // @[LoadQueue.scala 131:10:@4247.4]
  assign _T_3350 = 3'h5 <= offsetQ_0; // @[LoadQueue.scala 131:81:@4250.4]
  assign _T_3351 = _T_2848 & _T_3350; // @[LoadQueue.scala 131:72:@4251.4]
  assign _T_3353 = offsetQ_0 < 3'h5; // @[LoadQueue.scala 132:33:@4252.4]
  assign _T_3356 = _T_3353 & _T_2857; // @[LoadQueue.scala 132:41:@4254.4]
  assign _T_3358 = _T_3356 == 1'h0; // @[LoadQueue.scala 132:9:@4255.4]
  assign storesToCheck_0_5 = _T_1292 ? _T_3351 : _T_3358; // @[LoadQueue.scala 131:10:@4256.4]
  assign _T_3364 = 3'h6 <= offsetQ_0; // @[LoadQueue.scala 131:81:@4259.4]
  assign _T_3365 = _T_2865 & _T_3364; // @[LoadQueue.scala 131:72:@4260.4]
  assign _T_3367 = offsetQ_0 < 3'h6; // @[LoadQueue.scala 132:33:@4261.4]
  assign _T_3370 = _T_3367 & _T_2874; // @[LoadQueue.scala 132:41:@4263.4]
  assign _T_3372 = _T_3370 == 1'h0; // @[LoadQueue.scala 132:9:@4264.4]
  assign storesToCheck_0_6 = _T_1292 ? _T_3365 : _T_3372; // @[LoadQueue.scala 131:10:@4265.4]
  assign _T_3378 = 3'h7 <= offsetQ_0; // @[LoadQueue.scala 131:81:@4268.4]
  assign storesToCheck_0_7 = _T_1292 ? _T_3378 : 1'h1; // @[LoadQueue.scala 131:10:@4274.4]
  assign storesToCheck_1_0 = _T_1322 ? _T_2763 : 1'h1; // @[LoadQueue.scala 131:10:@4300.4]
  assign _T_3420 = 3'h1 <= offsetQ_1; // @[LoadQueue.scala 131:81:@4303.4]
  assign _T_3421 = _T_2780 & _T_3420; // @[LoadQueue.scala 131:72:@4304.4]
  assign _T_3423 = offsetQ_1 < 3'h1; // @[LoadQueue.scala 132:33:@4305.4]
  assign _T_3426 = _T_3423 & _T_2789; // @[LoadQueue.scala 132:41:@4307.4]
  assign _T_3428 = _T_3426 == 1'h0; // @[LoadQueue.scala 132:9:@4308.4]
  assign storesToCheck_1_1 = _T_1322 ? _T_3421 : _T_3428; // @[LoadQueue.scala 131:10:@4309.4]
  assign _T_3434 = 3'h2 <= offsetQ_1; // @[LoadQueue.scala 131:81:@4312.4]
  assign _T_3435 = _T_2797 & _T_3434; // @[LoadQueue.scala 131:72:@4313.4]
  assign _T_3437 = offsetQ_1 < 3'h2; // @[LoadQueue.scala 132:33:@4314.4]
  assign _T_3440 = _T_3437 & _T_2806; // @[LoadQueue.scala 132:41:@4316.4]
  assign _T_3442 = _T_3440 == 1'h0; // @[LoadQueue.scala 132:9:@4317.4]
  assign storesToCheck_1_2 = _T_1322 ? _T_3435 : _T_3442; // @[LoadQueue.scala 131:10:@4318.4]
  assign _T_3448 = 3'h3 <= offsetQ_1; // @[LoadQueue.scala 131:81:@4321.4]
  assign _T_3449 = _T_2814 & _T_3448; // @[LoadQueue.scala 131:72:@4322.4]
  assign _T_3451 = offsetQ_1 < 3'h3; // @[LoadQueue.scala 132:33:@4323.4]
  assign _T_3454 = _T_3451 & _T_2823; // @[LoadQueue.scala 132:41:@4325.4]
  assign _T_3456 = _T_3454 == 1'h0; // @[LoadQueue.scala 132:9:@4326.4]
  assign storesToCheck_1_3 = _T_1322 ? _T_3449 : _T_3456; // @[LoadQueue.scala 131:10:@4327.4]
  assign _T_3462 = 3'h4 <= offsetQ_1; // @[LoadQueue.scala 131:81:@4330.4]
  assign _T_3463 = _T_2831 & _T_3462; // @[LoadQueue.scala 131:72:@4331.4]
  assign _T_3465 = offsetQ_1 < 3'h4; // @[LoadQueue.scala 132:33:@4332.4]
  assign _T_3468 = _T_3465 & _T_2840; // @[LoadQueue.scala 132:41:@4334.4]
  assign _T_3470 = _T_3468 == 1'h0; // @[LoadQueue.scala 132:9:@4335.4]
  assign storesToCheck_1_4 = _T_1322 ? _T_3463 : _T_3470; // @[LoadQueue.scala 131:10:@4336.4]
  assign _T_3476 = 3'h5 <= offsetQ_1; // @[LoadQueue.scala 131:81:@4339.4]
  assign _T_3477 = _T_2848 & _T_3476; // @[LoadQueue.scala 131:72:@4340.4]
  assign _T_3479 = offsetQ_1 < 3'h5; // @[LoadQueue.scala 132:33:@4341.4]
  assign _T_3482 = _T_3479 & _T_2857; // @[LoadQueue.scala 132:41:@4343.4]
  assign _T_3484 = _T_3482 == 1'h0; // @[LoadQueue.scala 132:9:@4344.4]
  assign storesToCheck_1_5 = _T_1322 ? _T_3477 : _T_3484; // @[LoadQueue.scala 131:10:@4345.4]
  assign _T_3490 = 3'h6 <= offsetQ_1; // @[LoadQueue.scala 131:81:@4348.4]
  assign _T_3491 = _T_2865 & _T_3490; // @[LoadQueue.scala 131:72:@4349.4]
  assign _T_3493 = offsetQ_1 < 3'h6; // @[LoadQueue.scala 132:33:@4350.4]
  assign _T_3496 = _T_3493 & _T_2874; // @[LoadQueue.scala 132:41:@4352.4]
  assign _T_3498 = _T_3496 == 1'h0; // @[LoadQueue.scala 132:9:@4353.4]
  assign storesToCheck_1_6 = _T_1322 ? _T_3491 : _T_3498; // @[LoadQueue.scala 131:10:@4354.4]
  assign _T_3504 = 3'h7 <= offsetQ_1; // @[LoadQueue.scala 131:81:@4357.4]
  assign storesToCheck_1_7 = _T_1322 ? _T_3504 : 1'h1; // @[LoadQueue.scala 131:10:@4363.4]
  assign storesToCheck_2_0 = _T_1352 ? _T_2763 : 1'h1; // @[LoadQueue.scala 131:10:@4389.4]
  assign _T_3546 = 3'h1 <= offsetQ_2; // @[LoadQueue.scala 131:81:@4392.4]
  assign _T_3547 = _T_2780 & _T_3546; // @[LoadQueue.scala 131:72:@4393.4]
  assign _T_3549 = offsetQ_2 < 3'h1; // @[LoadQueue.scala 132:33:@4394.4]
  assign _T_3552 = _T_3549 & _T_2789; // @[LoadQueue.scala 132:41:@4396.4]
  assign _T_3554 = _T_3552 == 1'h0; // @[LoadQueue.scala 132:9:@4397.4]
  assign storesToCheck_2_1 = _T_1352 ? _T_3547 : _T_3554; // @[LoadQueue.scala 131:10:@4398.4]
  assign _T_3560 = 3'h2 <= offsetQ_2; // @[LoadQueue.scala 131:81:@4401.4]
  assign _T_3561 = _T_2797 & _T_3560; // @[LoadQueue.scala 131:72:@4402.4]
  assign _T_3563 = offsetQ_2 < 3'h2; // @[LoadQueue.scala 132:33:@4403.4]
  assign _T_3566 = _T_3563 & _T_2806; // @[LoadQueue.scala 132:41:@4405.4]
  assign _T_3568 = _T_3566 == 1'h0; // @[LoadQueue.scala 132:9:@4406.4]
  assign storesToCheck_2_2 = _T_1352 ? _T_3561 : _T_3568; // @[LoadQueue.scala 131:10:@4407.4]
  assign _T_3574 = 3'h3 <= offsetQ_2; // @[LoadQueue.scala 131:81:@4410.4]
  assign _T_3575 = _T_2814 & _T_3574; // @[LoadQueue.scala 131:72:@4411.4]
  assign _T_3577 = offsetQ_2 < 3'h3; // @[LoadQueue.scala 132:33:@4412.4]
  assign _T_3580 = _T_3577 & _T_2823; // @[LoadQueue.scala 132:41:@4414.4]
  assign _T_3582 = _T_3580 == 1'h0; // @[LoadQueue.scala 132:9:@4415.4]
  assign storesToCheck_2_3 = _T_1352 ? _T_3575 : _T_3582; // @[LoadQueue.scala 131:10:@4416.4]
  assign _T_3588 = 3'h4 <= offsetQ_2; // @[LoadQueue.scala 131:81:@4419.4]
  assign _T_3589 = _T_2831 & _T_3588; // @[LoadQueue.scala 131:72:@4420.4]
  assign _T_3591 = offsetQ_2 < 3'h4; // @[LoadQueue.scala 132:33:@4421.4]
  assign _T_3594 = _T_3591 & _T_2840; // @[LoadQueue.scala 132:41:@4423.4]
  assign _T_3596 = _T_3594 == 1'h0; // @[LoadQueue.scala 132:9:@4424.4]
  assign storesToCheck_2_4 = _T_1352 ? _T_3589 : _T_3596; // @[LoadQueue.scala 131:10:@4425.4]
  assign _T_3602 = 3'h5 <= offsetQ_2; // @[LoadQueue.scala 131:81:@4428.4]
  assign _T_3603 = _T_2848 & _T_3602; // @[LoadQueue.scala 131:72:@4429.4]
  assign _T_3605 = offsetQ_2 < 3'h5; // @[LoadQueue.scala 132:33:@4430.4]
  assign _T_3608 = _T_3605 & _T_2857; // @[LoadQueue.scala 132:41:@4432.4]
  assign _T_3610 = _T_3608 == 1'h0; // @[LoadQueue.scala 132:9:@4433.4]
  assign storesToCheck_2_5 = _T_1352 ? _T_3603 : _T_3610; // @[LoadQueue.scala 131:10:@4434.4]
  assign _T_3616 = 3'h6 <= offsetQ_2; // @[LoadQueue.scala 131:81:@4437.4]
  assign _T_3617 = _T_2865 & _T_3616; // @[LoadQueue.scala 131:72:@4438.4]
  assign _T_3619 = offsetQ_2 < 3'h6; // @[LoadQueue.scala 132:33:@4439.4]
  assign _T_3622 = _T_3619 & _T_2874; // @[LoadQueue.scala 132:41:@4441.4]
  assign _T_3624 = _T_3622 == 1'h0; // @[LoadQueue.scala 132:9:@4442.4]
  assign storesToCheck_2_6 = _T_1352 ? _T_3617 : _T_3624; // @[LoadQueue.scala 131:10:@4443.4]
  assign _T_3630 = 3'h7 <= offsetQ_2; // @[LoadQueue.scala 131:81:@4446.4]
  assign storesToCheck_2_7 = _T_1352 ? _T_3630 : 1'h1; // @[LoadQueue.scala 131:10:@4452.4]
  assign storesToCheck_3_0 = _T_1382 ? _T_2763 : 1'h1; // @[LoadQueue.scala 131:10:@4478.4]
  assign _T_3672 = 3'h1 <= offsetQ_3; // @[LoadQueue.scala 131:81:@4481.4]
  assign _T_3673 = _T_2780 & _T_3672; // @[LoadQueue.scala 131:72:@4482.4]
  assign _T_3675 = offsetQ_3 < 3'h1; // @[LoadQueue.scala 132:33:@4483.4]
  assign _T_3678 = _T_3675 & _T_2789; // @[LoadQueue.scala 132:41:@4485.4]
  assign _T_3680 = _T_3678 == 1'h0; // @[LoadQueue.scala 132:9:@4486.4]
  assign storesToCheck_3_1 = _T_1382 ? _T_3673 : _T_3680; // @[LoadQueue.scala 131:10:@4487.4]
  assign _T_3686 = 3'h2 <= offsetQ_3; // @[LoadQueue.scala 131:81:@4490.4]
  assign _T_3687 = _T_2797 & _T_3686; // @[LoadQueue.scala 131:72:@4491.4]
  assign _T_3689 = offsetQ_3 < 3'h2; // @[LoadQueue.scala 132:33:@4492.4]
  assign _T_3692 = _T_3689 & _T_2806; // @[LoadQueue.scala 132:41:@4494.4]
  assign _T_3694 = _T_3692 == 1'h0; // @[LoadQueue.scala 132:9:@4495.4]
  assign storesToCheck_3_2 = _T_1382 ? _T_3687 : _T_3694; // @[LoadQueue.scala 131:10:@4496.4]
  assign _T_3700 = 3'h3 <= offsetQ_3; // @[LoadQueue.scala 131:81:@4499.4]
  assign _T_3701 = _T_2814 & _T_3700; // @[LoadQueue.scala 131:72:@4500.4]
  assign _T_3703 = offsetQ_3 < 3'h3; // @[LoadQueue.scala 132:33:@4501.4]
  assign _T_3706 = _T_3703 & _T_2823; // @[LoadQueue.scala 132:41:@4503.4]
  assign _T_3708 = _T_3706 == 1'h0; // @[LoadQueue.scala 132:9:@4504.4]
  assign storesToCheck_3_3 = _T_1382 ? _T_3701 : _T_3708; // @[LoadQueue.scala 131:10:@4505.4]
  assign _T_3714 = 3'h4 <= offsetQ_3; // @[LoadQueue.scala 131:81:@4508.4]
  assign _T_3715 = _T_2831 & _T_3714; // @[LoadQueue.scala 131:72:@4509.4]
  assign _T_3717 = offsetQ_3 < 3'h4; // @[LoadQueue.scala 132:33:@4510.4]
  assign _T_3720 = _T_3717 & _T_2840; // @[LoadQueue.scala 132:41:@4512.4]
  assign _T_3722 = _T_3720 == 1'h0; // @[LoadQueue.scala 132:9:@4513.4]
  assign storesToCheck_3_4 = _T_1382 ? _T_3715 : _T_3722; // @[LoadQueue.scala 131:10:@4514.4]
  assign _T_3728 = 3'h5 <= offsetQ_3; // @[LoadQueue.scala 131:81:@4517.4]
  assign _T_3729 = _T_2848 & _T_3728; // @[LoadQueue.scala 131:72:@4518.4]
  assign _T_3731 = offsetQ_3 < 3'h5; // @[LoadQueue.scala 132:33:@4519.4]
  assign _T_3734 = _T_3731 & _T_2857; // @[LoadQueue.scala 132:41:@4521.4]
  assign _T_3736 = _T_3734 == 1'h0; // @[LoadQueue.scala 132:9:@4522.4]
  assign storesToCheck_3_5 = _T_1382 ? _T_3729 : _T_3736; // @[LoadQueue.scala 131:10:@4523.4]
  assign _T_3742 = 3'h6 <= offsetQ_3; // @[LoadQueue.scala 131:81:@4526.4]
  assign _T_3743 = _T_2865 & _T_3742; // @[LoadQueue.scala 131:72:@4527.4]
  assign _T_3745 = offsetQ_3 < 3'h6; // @[LoadQueue.scala 132:33:@4528.4]
  assign _T_3748 = _T_3745 & _T_2874; // @[LoadQueue.scala 132:41:@4530.4]
  assign _T_3750 = _T_3748 == 1'h0; // @[LoadQueue.scala 132:9:@4531.4]
  assign storesToCheck_3_6 = _T_1382 ? _T_3743 : _T_3750; // @[LoadQueue.scala 131:10:@4532.4]
  assign _T_3756 = 3'h7 <= offsetQ_3; // @[LoadQueue.scala 131:81:@4535.4]
  assign storesToCheck_3_7 = _T_1382 ? _T_3756 : 1'h1; // @[LoadQueue.scala 131:10:@4541.4]
  assign storesToCheck_4_0 = _T_1412 ? _T_2763 : 1'h1; // @[LoadQueue.scala 131:10:@4567.4]
  assign _T_3798 = 3'h1 <= offsetQ_4; // @[LoadQueue.scala 131:81:@4570.4]
  assign _T_3799 = _T_2780 & _T_3798; // @[LoadQueue.scala 131:72:@4571.4]
  assign _T_3801 = offsetQ_4 < 3'h1; // @[LoadQueue.scala 132:33:@4572.4]
  assign _T_3804 = _T_3801 & _T_2789; // @[LoadQueue.scala 132:41:@4574.4]
  assign _T_3806 = _T_3804 == 1'h0; // @[LoadQueue.scala 132:9:@4575.4]
  assign storesToCheck_4_1 = _T_1412 ? _T_3799 : _T_3806; // @[LoadQueue.scala 131:10:@4576.4]
  assign _T_3812 = 3'h2 <= offsetQ_4; // @[LoadQueue.scala 131:81:@4579.4]
  assign _T_3813 = _T_2797 & _T_3812; // @[LoadQueue.scala 131:72:@4580.4]
  assign _T_3815 = offsetQ_4 < 3'h2; // @[LoadQueue.scala 132:33:@4581.4]
  assign _T_3818 = _T_3815 & _T_2806; // @[LoadQueue.scala 132:41:@4583.4]
  assign _T_3820 = _T_3818 == 1'h0; // @[LoadQueue.scala 132:9:@4584.4]
  assign storesToCheck_4_2 = _T_1412 ? _T_3813 : _T_3820; // @[LoadQueue.scala 131:10:@4585.4]
  assign _T_3826 = 3'h3 <= offsetQ_4; // @[LoadQueue.scala 131:81:@4588.4]
  assign _T_3827 = _T_2814 & _T_3826; // @[LoadQueue.scala 131:72:@4589.4]
  assign _T_3829 = offsetQ_4 < 3'h3; // @[LoadQueue.scala 132:33:@4590.4]
  assign _T_3832 = _T_3829 & _T_2823; // @[LoadQueue.scala 132:41:@4592.4]
  assign _T_3834 = _T_3832 == 1'h0; // @[LoadQueue.scala 132:9:@4593.4]
  assign storesToCheck_4_3 = _T_1412 ? _T_3827 : _T_3834; // @[LoadQueue.scala 131:10:@4594.4]
  assign _T_3840 = 3'h4 <= offsetQ_4; // @[LoadQueue.scala 131:81:@4597.4]
  assign _T_3841 = _T_2831 & _T_3840; // @[LoadQueue.scala 131:72:@4598.4]
  assign _T_3843 = offsetQ_4 < 3'h4; // @[LoadQueue.scala 132:33:@4599.4]
  assign _T_3846 = _T_3843 & _T_2840; // @[LoadQueue.scala 132:41:@4601.4]
  assign _T_3848 = _T_3846 == 1'h0; // @[LoadQueue.scala 132:9:@4602.4]
  assign storesToCheck_4_4 = _T_1412 ? _T_3841 : _T_3848; // @[LoadQueue.scala 131:10:@4603.4]
  assign _T_3854 = 3'h5 <= offsetQ_4; // @[LoadQueue.scala 131:81:@4606.4]
  assign _T_3855 = _T_2848 & _T_3854; // @[LoadQueue.scala 131:72:@4607.4]
  assign _T_3857 = offsetQ_4 < 3'h5; // @[LoadQueue.scala 132:33:@4608.4]
  assign _T_3860 = _T_3857 & _T_2857; // @[LoadQueue.scala 132:41:@4610.4]
  assign _T_3862 = _T_3860 == 1'h0; // @[LoadQueue.scala 132:9:@4611.4]
  assign storesToCheck_4_5 = _T_1412 ? _T_3855 : _T_3862; // @[LoadQueue.scala 131:10:@4612.4]
  assign _T_3868 = 3'h6 <= offsetQ_4; // @[LoadQueue.scala 131:81:@4615.4]
  assign _T_3869 = _T_2865 & _T_3868; // @[LoadQueue.scala 131:72:@4616.4]
  assign _T_3871 = offsetQ_4 < 3'h6; // @[LoadQueue.scala 132:33:@4617.4]
  assign _T_3874 = _T_3871 & _T_2874; // @[LoadQueue.scala 132:41:@4619.4]
  assign _T_3876 = _T_3874 == 1'h0; // @[LoadQueue.scala 132:9:@4620.4]
  assign storesToCheck_4_6 = _T_1412 ? _T_3869 : _T_3876; // @[LoadQueue.scala 131:10:@4621.4]
  assign _T_3882 = 3'h7 <= offsetQ_4; // @[LoadQueue.scala 131:81:@4624.4]
  assign storesToCheck_4_7 = _T_1412 ? _T_3882 : 1'h1; // @[LoadQueue.scala 131:10:@4630.4]
  assign storesToCheck_5_0 = _T_1442 ? _T_2763 : 1'h1; // @[LoadQueue.scala 131:10:@4656.4]
  assign _T_3924 = 3'h1 <= offsetQ_5; // @[LoadQueue.scala 131:81:@4659.4]
  assign _T_3925 = _T_2780 & _T_3924; // @[LoadQueue.scala 131:72:@4660.4]
  assign _T_3927 = offsetQ_5 < 3'h1; // @[LoadQueue.scala 132:33:@4661.4]
  assign _T_3930 = _T_3927 & _T_2789; // @[LoadQueue.scala 132:41:@4663.4]
  assign _T_3932 = _T_3930 == 1'h0; // @[LoadQueue.scala 132:9:@4664.4]
  assign storesToCheck_5_1 = _T_1442 ? _T_3925 : _T_3932; // @[LoadQueue.scala 131:10:@4665.4]
  assign _T_3938 = 3'h2 <= offsetQ_5; // @[LoadQueue.scala 131:81:@4668.4]
  assign _T_3939 = _T_2797 & _T_3938; // @[LoadQueue.scala 131:72:@4669.4]
  assign _T_3941 = offsetQ_5 < 3'h2; // @[LoadQueue.scala 132:33:@4670.4]
  assign _T_3944 = _T_3941 & _T_2806; // @[LoadQueue.scala 132:41:@4672.4]
  assign _T_3946 = _T_3944 == 1'h0; // @[LoadQueue.scala 132:9:@4673.4]
  assign storesToCheck_5_2 = _T_1442 ? _T_3939 : _T_3946; // @[LoadQueue.scala 131:10:@4674.4]
  assign _T_3952 = 3'h3 <= offsetQ_5; // @[LoadQueue.scala 131:81:@4677.4]
  assign _T_3953 = _T_2814 & _T_3952; // @[LoadQueue.scala 131:72:@4678.4]
  assign _T_3955 = offsetQ_5 < 3'h3; // @[LoadQueue.scala 132:33:@4679.4]
  assign _T_3958 = _T_3955 & _T_2823; // @[LoadQueue.scala 132:41:@4681.4]
  assign _T_3960 = _T_3958 == 1'h0; // @[LoadQueue.scala 132:9:@4682.4]
  assign storesToCheck_5_3 = _T_1442 ? _T_3953 : _T_3960; // @[LoadQueue.scala 131:10:@4683.4]
  assign _T_3966 = 3'h4 <= offsetQ_5; // @[LoadQueue.scala 131:81:@4686.4]
  assign _T_3967 = _T_2831 & _T_3966; // @[LoadQueue.scala 131:72:@4687.4]
  assign _T_3969 = offsetQ_5 < 3'h4; // @[LoadQueue.scala 132:33:@4688.4]
  assign _T_3972 = _T_3969 & _T_2840; // @[LoadQueue.scala 132:41:@4690.4]
  assign _T_3974 = _T_3972 == 1'h0; // @[LoadQueue.scala 132:9:@4691.4]
  assign storesToCheck_5_4 = _T_1442 ? _T_3967 : _T_3974; // @[LoadQueue.scala 131:10:@4692.4]
  assign _T_3980 = 3'h5 <= offsetQ_5; // @[LoadQueue.scala 131:81:@4695.4]
  assign _T_3981 = _T_2848 & _T_3980; // @[LoadQueue.scala 131:72:@4696.4]
  assign _T_3983 = offsetQ_5 < 3'h5; // @[LoadQueue.scala 132:33:@4697.4]
  assign _T_3986 = _T_3983 & _T_2857; // @[LoadQueue.scala 132:41:@4699.4]
  assign _T_3988 = _T_3986 == 1'h0; // @[LoadQueue.scala 132:9:@4700.4]
  assign storesToCheck_5_5 = _T_1442 ? _T_3981 : _T_3988; // @[LoadQueue.scala 131:10:@4701.4]
  assign _T_3994 = 3'h6 <= offsetQ_5; // @[LoadQueue.scala 131:81:@4704.4]
  assign _T_3995 = _T_2865 & _T_3994; // @[LoadQueue.scala 131:72:@4705.4]
  assign _T_3997 = offsetQ_5 < 3'h6; // @[LoadQueue.scala 132:33:@4706.4]
  assign _T_4000 = _T_3997 & _T_2874; // @[LoadQueue.scala 132:41:@4708.4]
  assign _T_4002 = _T_4000 == 1'h0; // @[LoadQueue.scala 132:9:@4709.4]
  assign storesToCheck_5_6 = _T_1442 ? _T_3995 : _T_4002; // @[LoadQueue.scala 131:10:@4710.4]
  assign _T_4008 = 3'h7 <= offsetQ_5; // @[LoadQueue.scala 131:81:@4713.4]
  assign storesToCheck_5_7 = _T_1442 ? _T_4008 : 1'h1; // @[LoadQueue.scala 131:10:@4719.4]
  assign storesToCheck_6_0 = _T_1472 ? _T_2763 : 1'h1; // @[LoadQueue.scala 131:10:@4745.4]
  assign _T_4050 = 3'h1 <= offsetQ_6; // @[LoadQueue.scala 131:81:@4748.4]
  assign _T_4051 = _T_2780 & _T_4050; // @[LoadQueue.scala 131:72:@4749.4]
  assign _T_4053 = offsetQ_6 < 3'h1; // @[LoadQueue.scala 132:33:@4750.4]
  assign _T_4056 = _T_4053 & _T_2789; // @[LoadQueue.scala 132:41:@4752.4]
  assign _T_4058 = _T_4056 == 1'h0; // @[LoadQueue.scala 132:9:@4753.4]
  assign storesToCheck_6_1 = _T_1472 ? _T_4051 : _T_4058; // @[LoadQueue.scala 131:10:@4754.4]
  assign _T_4064 = 3'h2 <= offsetQ_6; // @[LoadQueue.scala 131:81:@4757.4]
  assign _T_4065 = _T_2797 & _T_4064; // @[LoadQueue.scala 131:72:@4758.4]
  assign _T_4067 = offsetQ_6 < 3'h2; // @[LoadQueue.scala 132:33:@4759.4]
  assign _T_4070 = _T_4067 & _T_2806; // @[LoadQueue.scala 132:41:@4761.4]
  assign _T_4072 = _T_4070 == 1'h0; // @[LoadQueue.scala 132:9:@4762.4]
  assign storesToCheck_6_2 = _T_1472 ? _T_4065 : _T_4072; // @[LoadQueue.scala 131:10:@4763.4]
  assign _T_4078 = 3'h3 <= offsetQ_6; // @[LoadQueue.scala 131:81:@4766.4]
  assign _T_4079 = _T_2814 & _T_4078; // @[LoadQueue.scala 131:72:@4767.4]
  assign _T_4081 = offsetQ_6 < 3'h3; // @[LoadQueue.scala 132:33:@4768.4]
  assign _T_4084 = _T_4081 & _T_2823; // @[LoadQueue.scala 132:41:@4770.4]
  assign _T_4086 = _T_4084 == 1'h0; // @[LoadQueue.scala 132:9:@4771.4]
  assign storesToCheck_6_3 = _T_1472 ? _T_4079 : _T_4086; // @[LoadQueue.scala 131:10:@4772.4]
  assign _T_4092 = 3'h4 <= offsetQ_6; // @[LoadQueue.scala 131:81:@4775.4]
  assign _T_4093 = _T_2831 & _T_4092; // @[LoadQueue.scala 131:72:@4776.4]
  assign _T_4095 = offsetQ_6 < 3'h4; // @[LoadQueue.scala 132:33:@4777.4]
  assign _T_4098 = _T_4095 & _T_2840; // @[LoadQueue.scala 132:41:@4779.4]
  assign _T_4100 = _T_4098 == 1'h0; // @[LoadQueue.scala 132:9:@4780.4]
  assign storesToCheck_6_4 = _T_1472 ? _T_4093 : _T_4100; // @[LoadQueue.scala 131:10:@4781.4]
  assign _T_4106 = 3'h5 <= offsetQ_6; // @[LoadQueue.scala 131:81:@4784.4]
  assign _T_4107 = _T_2848 & _T_4106; // @[LoadQueue.scala 131:72:@4785.4]
  assign _T_4109 = offsetQ_6 < 3'h5; // @[LoadQueue.scala 132:33:@4786.4]
  assign _T_4112 = _T_4109 & _T_2857; // @[LoadQueue.scala 132:41:@4788.4]
  assign _T_4114 = _T_4112 == 1'h0; // @[LoadQueue.scala 132:9:@4789.4]
  assign storesToCheck_6_5 = _T_1472 ? _T_4107 : _T_4114; // @[LoadQueue.scala 131:10:@4790.4]
  assign _T_4120 = 3'h6 <= offsetQ_6; // @[LoadQueue.scala 131:81:@4793.4]
  assign _T_4121 = _T_2865 & _T_4120; // @[LoadQueue.scala 131:72:@4794.4]
  assign _T_4123 = offsetQ_6 < 3'h6; // @[LoadQueue.scala 132:33:@4795.4]
  assign _T_4126 = _T_4123 & _T_2874; // @[LoadQueue.scala 132:41:@4797.4]
  assign _T_4128 = _T_4126 == 1'h0; // @[LoadQueue.scala 132:9:@4798.4]
  assign storesToCheck_6_6 = _T_1472 ? _T_4121 : _T_4128; // @[LoadQueue.scala 131:10:@4799.4]
  assign _T_4134 = 3'h7 <= offsetQ_6; // @[LoadQueue.scala 131:81:@4802.4]
  assign storesToCheck_6_7 = _T_1472 ? _T_4134 : 1'h1; // @[LoadQueue.scala 131:10:@4808.4]
  assign storesToCheck_7_0 = _T_1502 ? _T_2763 : 1'h1; // @[LoadQueue.scala 131:10:@4834.4]
  assign _T_4176 = 3'h1 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4837.4]
  assign _T_4177 = _T_2780 & _T_4176; // @[LoadQueue.scala 131:72:@4838.4]
  assign _T_4179 = offsetQ_7 < 3'h1; // @[LoadQueue.scala 132:33:@4839.4]
  assign _T_4182 = _T_4179 & _T_2789; // @[LoadQueue.scala 132:41:@4841.4]
  assign _T_4184 = _T_4182 == 1'h0; // @[LoadQueue.scala 132:9:@4842.4]
  assign storesToCheck_7_1 = _T_1502 ? _T_4177 : _T_4184; // @[LoadQueue.scala 131:10:@4843.4]
  assign _T_4190 = 3'h2 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4846.4]
  assign _T_4191 = _T_2797 & _T_4190; // @[LoadQueue.scala 131:72:@4847.4]
  assign _T_4193 = offsetQ_7 < 3'h2; // @[LoadQueue.scala 132:33:@4848.4]
  assign _T_4196 = _T_4193 & _T_2806; // @[LoadQueue.scala 132:41:@4850.4]
  assign _T_4198 = _T_4196 == 1'h0; // @[LoadQueue.scala 132:9:@4851.4]
  assign storesToCheck_7_2 = _T_1502 ? _T_4191 : _T_4198; // @[LoadQueue.scala 131:10:@4852.4]
  assign _T_4204 = 3'h3 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4855.4]
  assign _T_4205 = _T_2814 & _T_4204; // @[LoadQueue.scala 131:72:@4856.4]
  assign _T_4207 = offsetQ_7 < 3'h3; // @[LoadQueue.scala 132:33:@4857.4]
  assign _T_4210 = _T_4207 & _T_2823; // @[LoadQueue.scala 132:41:@4859.4]
  assign _T_4212 = _T_4210 == 1'h0; // @[LoadQueue.scala 132:9:@4860.4]
  assign storesToCheck_7_3 = _T_1502 ? _T_4205 : _T_4212; // @[LoadQueue.scala 131:10:@4861.4]
  assign _T_4218 = 3'h4 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4864.4]
  assign _T_4219 = _T_2831 & _T_4218; // @[LoadQueue.scala 131:72:@4865.4]
  assign _T_4221 = offsetQ_7 < 3'h4; // @[LoadQueue.scala 132:33:@4866.4]
  assign _T_4224 = _T_4221 & _T_2840; // @[LoadQueue.scala 132:41:@4868.4]
  assign _T_4226 = _T_4224 == 1'h0; // @[LoadQueue.scala 132:9:@4869.4]
  assign storesToCheck_7_4 = _T_1502 ? _T_4219 : _T_4226; // @[LoadQueue.scala 131:10:@4870.4]
  assign _T_4232 = 3'h5 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4873.4]
  assign _T_4233 = _T_2848 & _T_4232; // @[LoadQueue.scala 131:72:@4874.4]
  assign _T_4235 = offsetQ_7 < 3'h5; // @[LoadQueue.scala 132:33:@4875.4]
  assign _T_4238 = _T_4235 & _T_2857; // @[LoadQueue.scala 132:41:@4877.4]
  assign _T_4240 = _T_4238 == 1'h0; // @[LoadQueue.scala 132:9:@4878.4]
  assign storesToCheck_7_5 = _T_1502 ? _T_4233 : _T_4240; // @[LoadQueue.scala 131:10:@4879.4]
  assign _T_4246 = 3'h6 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4882.4]
  assign _T_4247 = _T_2865 & _T_4246; // @[LoadQueue.scala 131:72:@4883.4]
  assign _T_4249 = offsetQ_7 < 3'h6; // @[LoadQueue.scala 132:33:@4884.4]
  assign _T_4252 = _T_4249 & _T_2874; // @[LoadQueue.scala 132:41:@4886.4]
  assign _T_4254 = _T_4252 == 1'h0; // @[LoadQueue.scala 132:9:@4887.4]
  assign storesToCheck_7_6 = _T_1502 ? _T_4247 : _T_4254; // @[LoadQueue.scala 131:10:@4888.4]
  assign _T_4260 = 3'h7 <= offsetQ_7; // @[LoadQueue.scala 131:81:@4891.4]
  assign storesToCheck_7_7 = _T_1502 ? _T_4260 : 1'h1; // @[LoadQueue.scala 131:10:@4897.4]
  assign _T_4650 = storesToCheck_0_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4916.4]
  assign entriesToCheck_0_0 = _T_4650 & checkBits_0; // @[LoadQueue.scala 141:26:@4917.4]
  assign _T_4652 = storesToCheck_0_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4918.4]
  assign entriesToCheck_0_1 = _T_4652 & checkBits_0; // @[LoadQueue.scala 141:26:@4919.4]
  assign _T_4654 = storesToCheck_0_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4920.4]
  assign entriesToCheck_0_2 = _T_4654 & checkBits_0; // @[LoadQueue.scala 141:26:@4921.4]
  assign _T_4656 = storesToCheck_0_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4922.4]
  assign entriesToCheck_0_3 = _T_4656 & checkBits_0; // @[LoadQueue.scala 141:26:@4923.4]
  assign _T_4658 = storesToCheck_0_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4924.4]
  assign entriesToCheck_0_4 = _T_4658 & checkBits_0; // @[LoadQueue.scala 141:26:@4925.4]
  assign _T_4660 = storesToCheck_0_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4926.4]
  assign entriesToCheck_0_5 = _T_4660 & checkBits_0; // @[LoadQueue.scala 141:26:@4927.4]
  assign _T_4662 = storesToCheck_0_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4928.4]
  assign entriesToCheck_0_6 = _T_4662 & checkBits_0; // @[LoadQueue.scala 141:26:@4929.4]
  assign _T_4664 = storesToCheck_0_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4930.4]
  assign entriesToCheck_0_7 = _T_4664 & checkBits_0; // @[LoadQueue.scala 141:26:@4931.4]
  assign _T_4666 = storesToCheck_1_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4940.4]
  assign entriesToCheck_1_0 = _T_4666 & checkBits_1; // @[LoadQueue.scala 141:26:@4941.4]
  assign _T_4668 = storesToCheck_1_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4942.4]
  assign entriesToCheck_1_1 = _T_4668 & checkBits_1; // @[LoadQueue.scala 141:26:@4943.4]
  assign _T_4670 = storesToCheck_1_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4944.4]
  assign entriesToCheck_1_2 = _T_4670 & checkBits_1; // @[LoadQueue.scala 141:26:@4945.4]
  assign _T_4672 = storesToCheck_1_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4946.4]
  assign entriesToCheck_1_3 = _T_4672 & checkBits_1; // @[LoadQueue.scala 141:26:@4947.4]
  assign _T_4674 = storesToCheck_1_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4948.4]
  assign entriesToCheck_1_4 = _T_4674 & checkBits_1; // @[LoadQueue.scala 141:26:@4949.4]
  assign _T_4676 = storesToCheck_1_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4950.4]
  assign entriesToCheck_1_5 = _T_4676 & checkBits_1; // @[LoadQueue.scala 141:26:@4951.4]
  assign _T_4678 = storesToCheck_1_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4952.4]
  assign entriesToCheck_1_6 = _T_4678 & checkBits_1; // @[LoadQueue.scala 141:26:@4953.4]
  assign _T_4680 = storesToCheck_1_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4954.4]
  assign entriesToCheck_1_7 = _T_4680 & checkBits_1; // @[LoadQueue.scala 141:26:@4955.4]
  assign _T_4682 = storesToCheck_2_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4964.4]
  assign entriesToCheck_2_0 = _T_4682 & checkBits_2; // @[LoadQueue.scala 141:26:@4965.4]
  assign _T_4684 = storesToCheck_2_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4966.4]
  assign entriesToCheck_2_1 = _T_4684 & checkBits_2; // @[LoadQueue.scala 141:26:@4967.4]
  assign _T_4686 = storesToCheck_2_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4968.4]
  assign entriesToCheck_2_2 = _T_4686 & checkBits_2; // @[LoadQueue.scala 141:26:@4969.4]
  assign _T_4688 = storesToCheck_2_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4970.4]
  assign entriesToCheck_2_3 = _T_4688 & checkBits_2; // @[LoadQueue.scala 141:26:@4971.4]
  assign _T_4690 = storesToCheck_2_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4972.4]
  assign entriesToCheck_2_4 = _T_4690 & checkBits_2; // @[LoadQueue.scala 141:26:@4973.4]
  assign _T_4692 = storesToCheck_2_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4974.4]
  assign entriesToCheck_2_5 = _T_4692 & checkBits_2; // @[LoadQueue.scala 141:26:@4975.4]
  assign _T_4694 = storesToCheck_2_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@4976.4]
  assign entriesToCheck_2_6 = _T_4694 & checkBits_2; // @[LoadQueue.scala 141:26:@4977.4]
  assign _T_4696 = storesToCheck_2_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@4978.4]
  assign entriesToCheck_2_7 = _T_4696 & checkBits_2; // @[LoadQueue.scala 141:26:@4979.4]
  assign _T_4698 = storesToCheck_3_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@4988.4]
  assign entriesToCheck_3_0 = _T_4698 & checkBits_3; // @[LoadQueue.scala 141:26:@4989.4]
  assign _T_4700 = storesToCheck_3_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@4990.4]
  assign entriesToCheck_3_1 = _T_4700 & checkBits_3; // @[LoadQueue.scala 141:26:@4991.4]
  assign _T_4702 = storesToCheck_3_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@4992.4]
  assign entriesToCheck_3_2 = _T_4702 & checkBits_3; // @[LoadQueue.scala 141:26:@4993.4]
  assign _T_4704 = storesToCheck_3_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@4994.4]
  assign entriesToCheck_3_3 = _T_4704 & checkBits_3; // @[LoadQueue.scala 141:26:@4995.4]
  assign _T_4706 = storesToCheck_3_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@4996.4]
  assign entriesToCheck_3_4 = _T_4706 & checkBits_3; // @[LoadQueue.scala 141:26:@4997.4]
  assign _T_4708 = storesToCheck_3_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@4998.4]
  assign entriesToCheck_3_5 = _T_4708 & checkBits_3; // @[LoadQueue.scala 141:26:@4999.4]
  assign _T_4710 = storesToCheck_3_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@5000.4]
  assign entriesToCheck_3_6 = _T_4710 & checkBits_3; // @[LoadQueue.scala 141:26:@5001.4]
  assign _T_4712 = storesToCheck_3_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@5002.4]
  assign entriesToCheck_3_7 = _T_4712 & checkBits_3; // @[LoadQueue.scala 141:26:@5003.4]
  assign _T_4714 = storesToCheck_4_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@5012.4]
  assign entriesToCheck_4_0 = _T_4714 & checkBits_4; // @[LoadQueue.scala 141:26:@5013.4]
  assign _T_4716 = storesToCheck_4_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@5014.4]
  assign entriesToCheck_4_1 = _T_4716 & checkBits_4; // @[LoadQueue.scala 141:26:@5015.4]
  assign _T_4718 = storesToCheck_4_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@5016.4]
  assign entriesToCheck_4_2 = _T_4718 & checkBits_4; // @[LoadQueue.scala 141:26:@5017.4]
  assign _T_4720 = storesToCheck_4_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@5018.4]
  assign entriesToCheck_4_3 = _T_4720 & checkBits_4; // @[LoadQueue.scala 141:26:@5019.4]
  assign _T_4722 = storesToCheck_4_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@5020.4]
  assign entriesToCheck_4_4 = _T_4722 & checkBits_4; // @[LoadQueue.scala 141:26:@5021.4]
  assign _T_4724 = storesToCheck_4_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@5022.4]
  assign entriesToCheck_4_5 = _T_4724 & checkBits_4; // @[LoadQueue.scala 141:26:@5023.4]
  assign _T_4726 = storesToCheck_4_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@5024.4]
  assign entriesToCheck_4_6 = _T_4726 & checkBits_4; // @[LoadQueue.scala 141:26:@5025.4]
  assign _T_4728 = storesToCheck_4_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@5026.4]
  assign entriesToCheck_4_7 = _T_4728 & checkBits_4; // @[LoadQueue.scala 141:26:@5027.4]
  assign _T_4730 = storesToCheck_5_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@5036.4]
  assign entriesToCheck_5_0 = _T_4730 & checkBits_5; // @[LoadQueue.scala 141:26:@5037.4]
  assign _T_4732 = storesToCheck_5_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@5038.4]
  assign entriesToCheck_5_1 = _T_4732 & checkBits_5; // @[LoadQueue.scala 141:26:@5039.4]
  assign _T_4734 = storesToCheck_5_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@5040.4]
  assign entriesToCheck_5_2 = _T_4734 & checkBits_5; // @[LoadQueue.scala 141:26:@5041.4]
  assign _T_4736 = storesToCheck_5_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@5042.4]
  assign entriesToCheck_5_3 = _T_4736 & checkBits_5; // @[LoadQueue.scala 141:26:@5043.4]
  assign _T_4738 = storesToCheck_5_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@5044.4]
  assign entriesToCheck_5_4 = _T_4738 & checkBits_5; // @[LoadQueue.scala 141:26:@5045.4]
  assign _T_4740 = storesToCheck_5_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@5046.4]
  assign entriesToCheck_5_5 = _T_4740 & checkBits_5; // @[LoadQueue.scala 141:26:@5047.4]
  assign _T_4742 = storesToCheck_5_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@5048.4]
  assign entriesToCheck_5_6 = _T_4742 & checkBits_5; // @[LoadQueue.scala 141:26:@5049.4]
  assign _T_4744 = storesToCheck_5_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@5050.4]
  assign entriesToCheck_5_7 = _T_4744 & checkBits_5; // @[LoadQueue.scala 141:26:@5051.4]
  assign _T_4746 = storesToCheck_6_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@5060.4]
  assign entriesToCheck_6_0 = _T_4746 & checkBits_6; // @[LoadQueue.scala 141:26:@5061.4]
  assign _T_4748 = storesToCheck_6_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@5062.4]
  assign entriesToCheck_6_1 = _T_4748 & checkBits_6; // @[LoadQueue.scala 141:26:@5063.4]
  assign _T_4750 = storesToCheck_6_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@5064.4]
  assign entriesToCheck_6_2 = _T_4750 & checkBits_6; // @[LoadQueue.scala 141:26:@5065.4]
  assign _T_4752 = storesToCheck_6_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@5066.4]
  assign entriesToCheck_6_3 = _T_4752 & checkBits_6; // @[LoadQueue.scala 141:26:@5067.4]
  assign _T_4754 = storesToCheck_6_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@5068.4]
  assign entriesToCheck_6_4 = _T_4754 & checkBits_6; // @[LoadQueue.scala 141:26:@5069.4]
  assign _T_4756 = storesToCheck_6_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@5070.4]
  assign entriesToCheck_6_5 = _T_4756 & checkBits_6; // @[LoadQueue.scala 141:26:@5071.4]
  assign _T_4758 = storesToCheck_6_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@5072.4]
  assign entriesToCheck_6_6 = _T_4758 & checkBits_6; // @[LoadQueue.scala 141:26:@5073.4]
  assign _T_4760 = storesToCheck_6_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@5074.4]
  assign entriesToCheck_6_7 = _T_4760 & checkBits_6; // @[LoadQueue.scala 141:26:@5075.4]
  assign _T_4762 = storesToCheck_7_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@5084.4]
  assign entriesToCheck_7_0 = _T_4762 & checkBits_7; // @[LoadQueue.scala 141:26:@5085.4]
  assign _T_4764 = storesToCheck_7_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@5086.4]
  assign entriesToCheck_7_1 = _T_4764 & checkBits_7; // @[LoadQueue.scala 141:26:@5087.4]
  assign _T_4766 = storesToCheck_7_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@5088.4]
  assign entriesToCheck_7_2 = _T_4766 & checkBits_7; // @[LoadQueue.scala 141:26:@5089.4]
  assign _T_4768 = storesToCheck_7_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@5090.4]
  assign entriesToCheck_7_3 = _T_4768 & checkBits_7; // @[LoadQueue.scala 141:26:@5091.4]
  assign _T_4770 = storesToCheck_7_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@5092.4]
  assign entriesToCheck_7_4 = _T_4770 & checkBits_7; // @[LoadQueue.scala 141:26:@5093.4]
  assign _T_4772 = storesToCheck_7_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@5094.4]
  assign entriesToCheck_7_5 = _T_4772 & checkBits_7; // @[LoadQueue.scala 141:26:@5095.4]
  assign _T_4774 = storesToCheck_7_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@5096.4]
  assign entriesToCheck_7_6 = _T_4774 & checkBits_7; // @[LoadQueue.scala 141:26:@5097.4]
  assign _T_4776 = storesToCheck_7_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@5098.4]
  assign entriesToCheck_7_7 = _T_4776 & checkBits_7; // @[LoadQueue.scala 141:26:@5099.4]
  assign _T_5144 = entriesToCheck_0_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@5109.4]
  assign _T_5145 = _T_5144 & addrKnown_0; // @[LoadQueue.scala 152:41:@5110.4]
  assign _T_5146 = addrQ_0 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@5111.4]
  assign conflict_0_0 = _T_5145 & _T_5146; // @[LoadQueue.scala 152:68:@5112.4]
  assign _T_5148 = entriesToCheck_0_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@5114.4]
  assign _T_5149 = _T_5148 & addrKnown_0; // @[LoadQueue.scala 152:41:@5115.4]
  assign _T_5150 = addrQ_0 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@5116.4]
  assign conflict_0_1 = _T_5149 & _T_5150; // @[LoadQueue.scala 152:68:@5117.4]
  assign _T_5152 = entriesToCheck_0_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@5119.4]
  assign _T_5153 = _T_5152 & addrKnown_0; // @[LoadQueue.scala 152:41:@5120.4]
  assign _T_5154 = addrQ_0 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@5121.4]
  assign conflict_0_2 = _T_5153 & _T_5154; // @[LoadQueue.scala 152:68:@5122.4]
  assign _T_5156 = entriesToCheck_0_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@5124.4]
  assign _T_5157 = _T_5156 & addrKnown_0; // @[LoadQueue.scala 152:41:@5125.4]
  assign _T_5158 = addrQ_0 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@5126.4]
  assign conflict_0_3 = _T_5157 & _T_5158; // @[LoadQueue.scala 152:68:@5127.4]
  assign _T_5160 = entriesToCheck_0_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@5129.4]
  assign _T_5161 = _T_5160 & addrKnown_0; // @[LoadQueue.scala 152:41:@5130.4]
  assign _T_5162 = addrQ_0 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@5131.4]
  assign conflict_0_4 = _T_5161 & _T_5162; // @[LoadQueue.scala 152:68:@5132.4]
  assign _T_5164 = entriesToCheck_0_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@5134.4]
  assign _T_5165 = _T_5164 & addrKnown_0; // @[LoadQueue.scala 152:41:@5135.4]
  assign _T_5166 = addrQ_0 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@5136.4]
  assign conflict_0_5 = _T_5165 & _T_5166; // @[LoadQueue.scala 152:68:@5137.4]
  assign _T_5168 = entriesToCheck_0_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@5139.4]
  assign _T_5169 = _T_5168 & addrKnown_0; // @[LoadQueue.scala 152:41:@5140.4]
  assign _T_5170 = addrQ_0 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@5141.4]
  assign conflict_0_6 = _T_5169 & _T_5170; // @[LoadQueue.scala 152:68:@5142.4]
  assign _T_5172 = entriesToCheck_0_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@5144.4]
  assign _T_5173 = _T_5172 & addrKnown_0; // @[LoadQueue.scala 152:41:@5145.4]
  assign _T_5174 = addrQ_0 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@5146.4]
  assign conflict_0_7 = _T_5173 & _T_5174; // @[LoadQueue.scala 152:68:@5147.4]
  assign _T_5176 = entriesToCheck_1_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@5149.4]
  assign _T_5177 = _T_5176 & addrKnown_1; // @[LoadQueue.scala 152:41:@5150.4]
  assign _T_5178 = addrQ_1 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@5151.4]
  assign conflict_1_0 = _T_5177 & _T_5178; // @[LoadQueue.scala 152:68:@5152.4]
  assign _T_5180 = entriesToCheck_1_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@5154.4]
  assign _T_5181 = _T_5180 & addrKnown_1; // @[LoadQueue.scala 152:41:@5155.4]
  assign _T_5182 = addrQ_1 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@5156.4]
  assign conflict_1_1 = _T_5181 & _T_5182; // @[LoadQueue.scala 152:68:@5157.4]
  assign _T_5184 = entriesToCheck_1_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@5159.4]
  assign _T_5185 = _T_5184 & addrKnown_1; // @[LoadQueue.scala 152:41:@5160.4]
  assign _T_5186 = addrQ_1 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@5161.4]
  assign conflict_1_2 = _T_5185 & _T_5186; // @[LoadQueue.scala 152:68:@5162.4]
  assign _T_5188 = entriesToCheck_1_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@5164.4]
  assign _T_5189 = _T_5188 & addrKnown_1; // @[LoadQueue.scala 152:41:@5165.4]
  assign _T_5190 = addrQ_1 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@5166.4]
  assign conflict_1_3 = _T_5189 & _T_5190; // @[LoadQueue.scala 152:68:@5167.4]
  assign _T_5192 = entriesToCheck_1_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@5169.4]
  assign _T_5193 = _T_5192 & addrKnown_1; // @[LoadQueue.scala 152:41:@5170.4]
  assign _T_5194 = addrQ_1 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@5171.4]
  assign conflict_1_4 = _T_5193 & _T_5194; // @[LoadQueue.scala 152:68:@5172.4]
  assign _T_5196 = entriesToCheck_1_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@5174.4]
  assign _T_5197 = _T_5196 & addrKnown_1; // @[LoadQueue.scala 152:41:@5175.4]
  assign _T_5198 = addrQ_1 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@5176.4]
  assign conflict_1_5 = _T_5197 & _T_5198; // @[LoadQueue.scala 152:68:@5177.4]
  assign _T_5200 = entriesToCheck_1_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@5179.4]
  assign _T_5201 = _T_5200 & addrKnown_1; // @[LoadQueue.scala 152:41:@5180.4]
  assign _T_5202 = addrQ_1 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@5181.4]
  assign conflict_1_6 = _T_5201 & _T_5202; // @[LoadQueue.scala 152:68:@5182.4]
  assign _T_5204 = entriesToCheck_1_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@5184.4]
  assign _T_5205 = _T_5204 & addrKnown_1; // @[LoadQueue.scala 152:41:@5185.4]
  assign _T_5206 = addrQ_1 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@5186.4]
  assign conflict_1_7 = _T_5205 & _T_5206; // @[LoadQueue.scala 152:68:@5187.4]
  assign _T_5208 = entriesToCheck_2_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@5189.4]
  assign _T_5209 = _T_5208 & addrKnown_2; // @[LoadQueue.scala 152:41:@5190.4]
  assign _T_5210 = addrQ_2 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@5191.4]
  assign conflict_2_0 = _T_5209 & _T_5210; // @[LoadQueue.scala 152:68:@5192.4]
  assign _T_5212 = entriesToCheck_2_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@5194.4]
  assign _T_5213 = _T_5212 & addrKnown_2; // @[LoadQueue.scala 152:41:@5195.4]
  assign _T_5214 = addrQ_2 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@5196.4]
  assign conflict_2_1 = _T_5213 & _T_5214; // @[LoadQueue.scala 152:68:@5197.4]
  assign _T_5216 = entriesToCheck_2_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@5199.4]
  assign _T_5217 = _T_5216 & addrKnown_2; // @[LoadQueue.scala 152:41:@5200.4]
  assign _T_5218 = addrQ_2 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@5201.4]
  assign conflict_2_2 = _T_5217 & _T_5218; // @[LoadQueue.scala 152:68:@5202.4]
  assign _T_5220 = entriesToCheck_2_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@5204.4]
  assign _T_5221 = _T_5220 & addrKnown_2; // @[LoadQueue.scala 152:41:@5205.4]
  assign _T_5222 = addrQ_2 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@5206.4]
  assign conflict_2_3 = _T_5221 & _T_5222; // @[LoadQueue.scala 152:68:@5207.4]
  assign _T_5224 = entriesToCheck_2_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@5209.4]
  assign _T_5225 = _T_5224 & addrKnown_2; // @[LoadQueue.scala 152:41:@5210.4]
  assign _T_5226 = addrQ_2 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@5211.4]
  assign conflict_2_4 = _T_5225 & _T_5226; // @[LoadQueue.scala 152:68:@5212.4]
  assign _T_5228 = entriesToCheck_2_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@5214.4]
  assign _T_5229 = _T_5228 & addrKnown_2; // @[LoadQueue.scala 152:41:@5215.4]
  assign _T_5230 = addrQ_2 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@5216.4]
  assign conflict_2_5 = _T_5229 & _T_5230; // @[LoadQueue.scala 152:68:@5217.4]
  assign _T_5232 = entriesToCheck_2_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@5219.4]
  assign _T_5233 = _T_5232 & addrKnown_2; // @[LoadQueue.scala 152:41:@5220.4]
  assign _T_5234 = addrQ_2 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@5221.4]
  assign conflict_2_6 = _T_5233 & _T_5234; // @[LoadQueue.scala 152:68:@5222.4]
  assign _T_5236 = entriesToCheck_2_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@5224.4]
  assign _T_5237 = _T_5236 & addrKnown_2; // @[LoadQueue.scala 152:41:@5225.4]
  assign _T_5238 = addrQ_2 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@5226.4]
  assign conflict_2_7 = _T_5237 & _T_5238; // @[LoadQueue.scala 152:68:@5227.4]
  assign _T_5240 = entriesToCheck_3_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@5229.4]
  assign _T_5241 = _T_5240 & addrKnown_3; // @[LoadQueue.scala 152:41:@5230.4]
  assign _T_5242 = addrQ_3 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@5231.4]
  assign conflict_3_0 = _T_5241 & _T_5242; // @[LoadQueue.scala 152:68:@5232.4]
  assign _T_5244 = entriesToCheck_3_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@5234.4]
  assign _T_5245 = _T_5244 & addrKnown_3; // @[LoadQueue.scala 152:41:@5235.4]
  assign _T_5246 = addrQ_3 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@5236.4]
  assign conflict_3_1 = _T_5245 & _T_5246; // @[LoadQueue.scala 152:68:@5237.4]
  assign _T_5248 = entriesToCheck_3_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@5239.4]
  assign _T_5249 = _T_5248 & addrKnown_3; // @[LoadQueue.scala 152:41:@5240.4]
  assign _T_5250 = addrQ_3 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@5241.4]
  assign conflict_3_2 = _T_5249 & _T_5250; // @[LoadQueue.scala 152:68:@5242.4]
  assign _T_5252 = entriesToCheck_3_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@5244.4]
  assign _T_5253 = _T_5252 & addrKnown_3; // @[LoadQueue.scala 152:41:@5245.4]
  assign _T_5254 = addrQ_3 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@5246.4]
  assign conflict_3_3 = _T_5253 & _T_5254; // @[LoadQueue.scala 152:68:@5247.4]
  assign _T_5256 = entriesToCheck_3_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@5249.4]
  assign _T_5257 = _T_5256 & addrKnown_3; // @[LoadQueue.scala 152:41:@5250.4]
  assign _T_5258 = addrQ_3 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@5251.4]
  assign conflict_3_4 = _T_5257 & _T_5258; // @[LoadQueue.scala 152:68:@5252.4]
  assign _T_5260 = entriesToCheck_3_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@5254.4]
  assign _T_5261 = _T_5260 & addrKnown_3; // @[LoadQueue.scala 152:41:@5255.4]
  assign _T_5262 = addrQ_3 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@5256.4]
  assign conflict_3_5 = _T_5261 & _T_5262; // @[LoadQueue.scala 152:68:@5257.4]
  assign _T_5264 = entriesToCheck_3_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@5259.4]
  assign _T_5265 = _T_5264 & addrKnown_3; // @[LoadQueue.scala 152:41:@5260.4]
  assign _T_5266 = addrQ_3 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@5261.4]
  assign conflict_3_6 = _T_5265 & _T_5266; // @[LoadQueue.scala 152:68:@5262.4]
  assign _T_5268 = entriesToCheck_3_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@5264.4]
  assign _T_5269 = _T_5268 & addrKnown_3; // @[LoadQueue.scala 152:41:@5265.4]
  assign _T_5270 = addrQ_3 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@5266.4]
  assign conflict_3_7 = _T_5269 & _T_5270; // @[LoadQueue.scala 152:68:@5267.4]
  assign _T_5272 = entriesToCheck_4_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@5269.4]
  assign _T_5273 = _T_5272 & addrKnown_4; // @[LoadQueue.scala 152:41:@5270.4]
  assign _T_5274 = addrQ_4 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@5271.4]
  assign conflict_4_0 = _T_5273 & _T_5274; // @[LoadQueue.scala 152:68:@5272.4]
  assign _T_5276 = entriesToCheck_4_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@5274.4]
  assign _T_5277 = _T_5276 & addrKnown_4; // @[LoadQueue.scala 152:41:@5275.4]
  assign _T_5278 = addrQ_4 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@5276.4]
  assign conflict_4_1 = _T_5277 & _T_5278; // @[LoadQueue.scala 152:68:@5277.4]
  assign _T_5280 = entriesToCheck_4_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@5279.4]
  assign _T_5281 = _T_5280 & addrKnown_4; // @[LoadQueue.scala 152:41:@5280.4]
  assign _T_5282 = addrQ_4 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@5281.4]
  assign conflict_4_2 = _T_5281 & _T_5282; // @[LoadQueue.scala 152:68:@5282.4]
  assign _T_5284 = entriesToCheck_4_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@5284.4]
  assign _T_5285 = _T_5284 & addrKnown_4; // @[LoadQueue.scala 152:41:@5285.4]
  assign _T_5286 = addrQ_4 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@5286.4]
  assign conflict_4_3 = _T_5285 & _T_5286; // @[LoadQueue.scala 152:68:@5287.4]
  assign _T_5288 = entriesToCheck_4_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@5289.4]
  assign _T_5289 = _T_5288 & addrKnown_4; // @[LoadQueue.scala 152:41:@5290.4]
  assign _T_5290 = addrQ_4 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@5291.4]
  assign conflict_4_4 = _T_5289 & _T_5290; // @[LoadQueue.scala 152:68:@5292.4]
  assign _T_5292 = entriesToCheck_4_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@5294.4]
  assign _T_5293 = _T_5292 & addrKnown_4; // @[LoadQueue.scala 152:41:@5295.4]
  assign _T_5294 = addrQ_4 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@5296.4]
  assign conflict_4_5 = _T_5293 & _T_5294; // @[LoadQueue.scala 152:68:@5297.4]
  assign _T_5296 = entriesToCheck_4_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@5299.4]
  assign _T_5297 = _T_5296 & addrKnown_4; // @[LoadQueue.scala 152:41:@5300.4]
  assign _T_5298 = addrQ_4 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@5301.4]
  assign conflict_4_6 = _T_5297 & _T_5298; // @[LoadQueue.scala 152:68:@5302.4]
  assign _T_5300 = entriesToCheck_4_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@5304.4]
  assign _T_5301 = _T_5300 & addrKnown_4; // @[LoadQueue.scala 152:41:@5305.4]
  assign _T_5302 = addrQ_4 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@5306.4]
  assign conflict_4_7 = _T_5301 & _T_5302; // @[LoadQueue.scala 152:68:@5307.4]
  assign _T_5304 = entriesToCheck_5_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@5309.4]
  assign _T_5305 = _T_5304 & addrKnown_5; // @[LoadQueue.scala 152:41:@5310.4]
  assign _T_5306 = addrQ_5 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@5311.4]
  assign conflict_5_0 = _T_5305 & _T_5306; // @[LoadQueue.scala 152:68:@5312.4]
  assign _T_5308 = entriesToCheck_5_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@5314.4]
  assign _T_5309 = _T_5308 & addrKnown_5; // @[LoadQueue.scala 152:41:@5315.4]
  assign _T_5310 = addrQ_5 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@5316.4]
  assign conflict_5_1 = _T_5309 & _T_5310; // @[LoadQueue.scala 152:68:@5317.4]
  assign _T_5312 = entriesToCheck_5_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@5319.4]
  assign _T_5313 = _T_5312 & addrKnown_5; // @[LoadQueue.scala 152:41:@5320.4]
  assign _T_5314 = addrQ_5 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@5321.4]
  assign conflict_5_2 = _T_5313 & _T_5314; // @[LoadQueue.scala 152:68:@5322.4]
  assign _T_5316 = entriesToCheck_5_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@5324.4]
  assign _T_5317 = _T_5316 & addrKnown_5; // @[LoadQueue.scala 152:41:@5325.4]
  assign _T_5318 = addrQ_5 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@5326.4]
  assign conflict_5_3 = _T_5317 & _T_5318; // @[LoadQueue.scala 152:68:@5327.4]
  assign _T_5320 = entriesToCheck_5_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@5329.4]
  assign _T_5321 = _T_5320 & addrKnown_5; // @[LoadQueue.scala 152:41:@5330.4]
  assign _T_5322 = addrQ_5 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@5331.4]
  assign conflict_5_4 = _T_5321 & _T_5322; // @[LoadQueue.scala 152:68:@5332.4]
  assign _T_5324 = entriesToCheck_5_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@5334.4]
  assign _T_5325 = _T_5324 & addrKnown_5; // @[LoadQueue.scala 152:41:@5335.4]
  assign _T_5326 = addrQ_5 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@5336.4]
  assign conflict_5_5 = _T_5325 & _T_5326; // @[LoadQueue.scala 152:68:@5337.4]
  assign _T_5328 = entriesToCheck_5_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@5339.4]
  assign _T_5329 = _T_5328 & addrKnown_5; // @[LoadQueue.scala 152:41:@5340.4]
  assign _T_5330 = addrQ_5 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@5341.4]
  assign conflict_5_6 = _T_5329 & _T_5330; // @[LoadQueue.scala 152:68:@5342.4]
  assign _T_5332 = entriesToCheck_5_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@5344.4]
  assign _T_5333 = _T_5332 & addrKnown_5; // @[LoadQueue.scala 152:41:@5345.4]
  assign _T_5334 = addrQ_5 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@5346.4]
  assign conflict_5_7 = _T_5333 & _T_5334; // @[LoadQueue.scala 152:68:@5347.4]
  assign _T_5336 = entriesToCheck_6_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@5349.4]
  assign _T_5337 = _T_5336 & addrKnown_6; // @[LoadQueue.scala 152:41:@5350.4]
  assign _T_5338 = addrQ_6 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@5351.4]
  assign conflict_6_0 = _T_5337 & _T_5338; // @[LoadQueue.scala 152:68:@5352.4]
  assign _T_5340 = entriesToCheck_6_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@5354.4]
  assign _T_5341 = _T_5340 & addrKnown_6; // @[LoadQueue.scala 152:41:@5355.4]
  assign _T_5342 = addrQ_6 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@5356.4]
  assign conflict_6_1 = _T_5341 & _T_5342; // @[LoadQueue.scala 152:68:@5357.4]
  assign _T_5344 = entriesToCheck_6_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@5359.4]
  assign _T_5345 = _T_5344 & addrKnown_6; // @[LoadQueue.scala 152:41:@5360.4]
  assign _T_5346 = addrQ_6 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@5361.4]
  assign conflict_6_2 = _T_5345 & _T_5346; // @[LoadQueue.scala 152:68:@5362.4]
  assign _T_5348 = entriesToCheck_6_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@5364.4]
  assign _T_5349 = _T_5348 & addrKnown_6; // @[LoadQueue.scala 152:41:@5365.4]
  assign _T_5350 = addrQ_6 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@5366.4]
  assign conflict_6_3 = _T_5349 & _T_5350; // @[LoadQueue.scala 152:68:@5367.4]
  assign _T_5352 = entriesToCheck_6_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@5369.4]
  assign _T_5353 = _T_5352 & addrKnown_6; // @[LoadQueue.scala 152:41:@5370.4]
  assign _T_5354 = addrQ_6 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@5371.4]
  assign conflict_6_4 = _T_5353 & _T_5354; // @[LoadQueue.scala 152:68:@5372.4]
  assign _T_5356 = entriesToCheck_6_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@5374.4]
  assign _T_5357 = _T_5356 & addrKnown_6; // @[LoadQueue.scala 152:41:@5375.4]
  assign _T_5358 = addrQ_6 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@5376.4]
  assign conflict_6_5 = _T_5357 & _T_5358; // @[LoadQueue.scala 152:68:@5377.4]
  assign _T_5360 = entriesToCheck_6_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@5379.4]
  assign _T_5361 = _T_5360 & addrKnown_6; // @[LoadQueue.scala 152:41:@5380.4]
  assign _T_5362 = addrQ_6 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@5381.4]
  assign conflict_6_6 = _T_5361 & _T_5362; // @[LoadQueue.scala 152:68:@5382.4]
  assign _T_5364 = entriesToCheck_6_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@5384.4]
  assign _T_5365 = _T_5364 & addrKnown_6; // @[LoadQueue.scala 152:41:@5385.4]
  assign _T_5366 = addrQ_6 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@5386.4]
  assign conflict_6_7 = _T_5365 & _T_5366; // @[LoadQueue.scala 152:68:@5387.4]
  assign _T_5368 = entriesToCheck_7_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@5389.4]
  assign _T_5369 = _T_5368 & addrKnown_7; // @[LoadQueue.scala 152:41:@5390.4]
  assign _T_5370 = addrQ_7 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@5391.4]
  assign conflict_7_0 = _T_5369 & _T_5370; // @[LoadQueue.scala 152:68:@5392.4]
  assign _T_5372 = entriesToCheck_7_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@5394.4]
  assign _T_5373 = _T_5372 & addrKnown_7; // @[LoadQueue.scala 152:41:@5395.4]
  assign _T_5374 = addrQ_7 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@5396.4]
  assign conflict_7_1 = _T_5373 & _T_5374; // @[LoadQueue.scala 152:68:@5397.4]
  assign _T_5376 = entriesToCheck_7_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@5399.4]
  assign _T_5377 = _T_5376 & addrKnown_7; // @[LoadQueue.scala 152:41:@5400.4]
  assign _T_5378 = addrQ_7 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@5401.4]
  assign conflict_7_2 = _T_5377 & _T_5378; // @[LoadQueue.scala 152:68:@5402.4]
  assign _T_5380 = entriesToCheck_7_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@5404.4]
  assign _T_5381 = _T_5380 & addrKnown_7; // @[LoadQueue.scala 152:41:@5405.4]
  assign _T_5382 = addrQ_7 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@5406.4]
  assign conflict_7_3 = _T_5381 & _T_5382; // @[LoadQueue.scala 152:68:@5407.4]
  assign _T_5384 = entriesToCheck_7_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@5409.4]
  assign _T_5385 = _T_5384 & addrKnown_7; // @[LoadQueue.scala 152:41:@5410.4]
  assign _T_5386 = addrQ_7 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@5411.4]
  assign conflict_7_4 = _T_5385 & _T_5386; // @[LoadQueue.scala 152:68:@5412.4]
  assign _T_5388 = entriesToCheck_7_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@5414.4]
  assign _T_5389 = _T_5388 & addrKnown_7; // @[LoadQueue.scala 152:41:@5415.4]
  assign _T_5390 = addrQ_7 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@5416.4]
  assign conflict_7_5 = _T_5389 & _T_5390; // @[LoadQueue.scala 152:68:@5417.4]
  assign _T_5392 = entriesToCheck_7_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@5419.4]
  assign _T_5393 = _T_5392 & addrKnown_7; // @[LoadQueue.scala 152:41:@5420.4]
  assign _T_5394 = addrQ_7 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@5421.4]
  assign conflict_7_6 = _T_5393 & _T_5394; // @[LoadQueue.scala 152:68:@5422.4]
  assign _T_5396 = entriesToCheck_7_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@5424.4]
  assign _T_5397 = _T_5396 & addrKnown_7; // @[LoadQueue.scala 152:41:@5425.4]
  assign _T_5398 = addrQ_7 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@5426.4]
  assign conflict_7_7 = _T_5397 & _T_5398; // @[LoadQueue.scala 152:68:@5427.4]
  assign _T_5767 = io_storeAddrDone_0 == 1'h0; // @[LoadQueue.scala 163:13:@5430.4]
  assign storeAddrNotKnownFlags_0_0 = _T_5767 & entriesToCheck_0_0; // @[LoadQueue.scala 163:19:@5431.4]
  assign _T_5770 = io_storeAddrDone_1 == 1'h0; // @[LoadQueue.scala 163:13:@5432.4]
  assign storeAddrNotKnownFlags_0_1 = _T_5770 & entriesToCheck_0_1; // @[LoadQueue.scala 163:19:@5433.4]
  assign _T_5773 = io_storeAddrDone_2 == 1'h0; // @[LoadQueue.scala 163:13:@5434.4]
  assign storeAddrNotKnownFlags_0_2 = _T_5773 & entriesToCheck_0_2; // @[LoadQueue.scala 163:19:@5435.4]
  assign _T_5776 = io_storeAddrDone_3 == 1'h0; // @[LoadQueue.scala 163:13:@5436.4]
  assign storeAddrNotKnownFlags_0_3 = _T_5776 & entriesToCheck_0_3; // @[LoadQueue.scala 163:19:@5437.4]
  assign _T_5779 = io_storeAddrDone_4 == 1'h0; // @[LoadQueue.scala 163:13:@5438.4]
  assign storeAddrNotKnownFlags_0_4 = _T_5779 & entriesToCheck_0_4; // @[LoadQueue.scala 163:19:@5439.4]
  assign _T_5782 = io_storeAddrDone_5 == 1'h0; // @[LoadQueue.scala 163:13:@5440.4]
  assign storeAddrNotKnownFlags_0_5 = _T_5782 & entriesToCheck_0_5; // @[LoadQueue.scala 163:19:@5441.4]
  assign _T_5785 = io_storeAddrDone_6 == 1'h0; // @[LoadQueue.scala 163:13:@5442.4]
  assign storeAddrNotKnownFlags_0_6 = _T_5785 & entriesToCheck_0_6; // @[LoadQueue.scala 163:19:@5443.4]
  assign _T_5788 = io_storeAddrDone_7 == 1'h0; // @[LoadQueue.scala 163:13:@5444.4]
  assign storeAddrNotKnownFlags_0_7 = _T_5788 & entriesToCheck_0_7; // @[LoadQueue.scala 163:19:@5445.4]
  assign storeAddrNotKnownFlags_1_0 = _T_5767 & entriesToCheck_1_0; // @[LoadQueue.scala 163:19:@5455.4]
  assign storeAddrNotKnownFlags_1_1 = _T_5770 & entriesToCheck_1_1; // @[LoadQueue.scala 163:19:@5457.4]
  assign storeAddrNotKnownFlags_1_2 = _T_5773 & entriesToCheck_1_2; // @[LoadQueue.scala 163:19:@5459.4]
  assign storeAddrNotKnownFlags_1_3 = _T_5776 & entriesToCheck_1_3; // @[LoadQueue.scala 163:19:@5461.4]
  assign storeAddrNotKnownFlags_1_4 = _T_5779 & entriesToCheck_1_4; // @[LoadQueue.scala 163:19:@5463.4]
  assign storeAddrNotKnownFlags_1_5 = _T_5782 & entriesToCheck_1_5; // @[LoadQueue.scala 163:19:@5465.4]
  assign storeAddrNotKnownFlags_1_6 = _T_5785 & entriesToCheck_1_6; // @[LoadQueue.scala 163:19:@5467.4]
  assign storeAddrNotKnownFlags_1_7 = _T_5788 & entriesToCheck_1_7; // @[LoadQueue.scala 163:19:@5469.4]
  assign storeAddrNotKnownFlags_2_0 = _T_5767 & entriesToCheck_2_0; // @[LoadQueue.scala 163:19:@5479.4]
  assign storeAddrNotKnownFlags_2_1 = _T_5770 & entriesToCheck_2_1; // @[LoadQueue.scala 163:19:@5481.4]
  assign storeAddrNotKnownFlags_2_2 = _T_5773 & entriesToCheck_2_2; // @[LoadQueue.scala 163:19:@5483.4]
  assign storeAddrNotKnownFlags_2_3 = _T_5776 & entriesToCheck_2_3; // @[LoadQueue.scala 163:19:@5485.4]
  assign storeAddrNotKnownFlags_2_4 = _T_5779 & entriesToCheck_2_4; // @[LoadQueue.scala 163:19:@5487.4]
  assign storeAddrNotKnownFlags_2_5 = _T_5782 & entriesToCheck_2_5; // @[LoadQueue.scala 163:19:@5489.4]
  assign storeAddrNotKnownFlags_2_6 = _T_5785 & entriesToCheck_2_6; // @[LoadQueue.scala 163:19:@5491.4]
  assign storeAddrNotKnownFlags_2_7 = _T_5788 & entriesToCheck_2_7; // @[LoadQueue.scala 163:19:@5493.4]
  assign storeAddrNotKnownFlags_3_0 = _T_5767 & entriesToCheck_3_0; // @[LoadQueue.scala 163:19:@5503.4]
  assign storeAddrNotKnownFlags_3_1 = _T_5770 & entriesToCheck_3_1; // @[LoadQueue.scala 163:19:@5505.4]
  assign storeAddrNotKnownFlags_3_2 = _T_5773 & entriesToCheck_3_2; // @[LoadQueue.scala 163:19:@5507.4]
  assign storeAddrNotKnownFlags_3_3 = _T_5776 & entriesToCheck_3_3; // @[LoadQueue.scala 163:19:@5509.4]
  assign storeAddrNotKnownFlags_3_4 = _T_5779 & entriesToCheck_3_4; // @[LoadQueue.scala 163:19:@5511.4]
  assign storeAddrNotKnownFlags_3_5 = _T_5782 & entriesToCheck_3_5; // @[LoadQueue.scala 163:19:@5513.4]
  assign storeAddrNotKnownFlags_3_6 = _T_5785 & entriesToCheck_3_6; // @[LoadQueue.scala 163:19:@5515.4]
  assign storeAddrNotKnownFlags_3_7 = _T_5788 & entriesToCheck_3_7; // @[LoadQueue.scala 163:19:@5517.4]
  assign storeAddrNotKnownFlags_4_0 = _T_5767 & entriesToCheck_4_0; // @[LoadQueue.scala 163:19:@5527.4]
  assign storeAddrNotKnownFlags_4_1 = _T_5770 & entriesToCheck_4_1; // @[LoadQueue.scala 163:19:@5529.4]
  assign storeAddrNotKnownFlags_4_2 = _T_5773 & entriesToCheck_4_2; // @[LoadQueue.scala 163:19:@5531.4]
  assign storeAddrNotKnownFlags_4_3 = _T_5776 & entriesToCheck_4_3; // @[LoadQueue.scala 163:19:@5533.4]
  assign storeAddrNotKnownFlags_4_4 = _T_5779 & entriesToCheck_4_4; // @[LoadQueue.scala 163:19:@5535.4]
  assign storeAddrNotKnownFlags_4_5 = _T_5782 & entriesToCheck_4_5; // @[LoadQueue.scala 163:19:@5537.4]
  assign storeAddrNotKnownFlags_4_6 = _T_5785 & entriesToCheck_4_6; // @[LoadQueue.scala 163:19:@5539.4]
  assign storeAddrNotKnownFlags_4_7 = _T_5788 & entriesToCheck_4_7; // @[LoadQueue.scala 163:19:@5541.4]
  assign storeAddrNotKnownFlags_5_0 = _T_5767 & entriesToCheck_5_0; // @[LoadQueue.scala 163:19:@5551.4]
  assign storeAddrNotKnownFlags_5_1 = _T_5770 & entriesToCheck_5_1; // @[LoadQueue.scala 163:19:@5553.4]
  assign storeAddrNotKnownFlags_5_2 = _T_5773 & entriesToCheck_5_2; // @[LoadQueue.scala 163:19:@5555.4]
  assign storeAddrNotKnownFlags_5_3 = _T_5776 & entriesToCheck_5_3; // @[LoadQueue.scala 163:19:@5557.4]
  assign storeAddrNotKnownFlags_5_4 = _T_5779 & entriesToCheck_5_4; // @[LoadQueue.scala 163:19:@5559.4]
  assign storeAddrNotKnownFlags_5_5 = _T_5782 & entriesToCheck_5_5; // @[LoadQueue.scala 163:19:@5561.4]
  assign storeAddrNotKnownFlags_5_6 = _T_5785 & entriesToCheck_5_6; // @[LoadQueue.scala 163:19:@5563.4]
  assign storeAddrNotKnownFlags_5_7 = _T_5788 & entriesToCheck_5_7; // @[LoadQueue.scala 163:19:@5565.4]
  assign storeAddrNotKnownFlags_6_0 = _T_5767 & entriesToCheck_6_0; // @[LoadQueue.scala 163:19:@5575.4]
  assign storeAddrNotKnownFlags_6_1 = _T_5770 & entriesToCheck_6_1; // @[LoadQueue.scala 163:19:@5577.4]
  assign storeAddrNotKnownFlags_6_2 = _T_5773 & entriesToCheck_6_2; // @[LoadQueue.scala 163:19:@5579.4]
  assign storeAddrNotKnownFlags_6_3 = _T_5776 & entriesToCheck_6_3; // @[LoadQueue.scala 163:19:@5581.4]
  assign storeAddrNotKnownFlags_6_4 = _T_5779 & entriesToCheck_6_4; // @[LoadQueue.scala 163:19:@5583.4]
  assign storeAddrNotKnownFlags_6_5 = _T_5782 & entriesToCheck_6_5; // @[LoadQueue.scala 163:19:@5585.4]
  assign storeAddrNotKnownFlags_6_6 = _T_5785 & entriesToCheck_6_6; // @[LoadQueue.scala 163:19:@5587.4]
  assign storeAddrNotKnownFlags_6_7 = _T_5788 & entriesToCheck_6_7; // @[LoadQueue.scala 163:19:@5589.4]
  assign storeAddrNotKnownFlags_7_0 = _T_5767 & entriesToCheck_7_0; // @[LoadQueue.scala 163:19:@5599.4]
  assign storeAddrNotKnownFlags_7_1 = _T_5770 & entriesToCheck_7_1; // @[LoadQueue.scala 163:19:@5601.4]
  assign storeAddrNotKnownFlags_7_2 = _T_5773 & entriesToCheck_7_2; // @[LoadQueue.scala 163:19:@5603.4]
  assign storeAddrNotKnownFlags_7_3 = _T_5776 & entriesToCheck_7_3; // @[LoadQueue.scala 163:19:@5605.4]
  assign storeAddrNotKnownFlags_7_4 = _T_5779 & entriesToCheck_7_4; // @[LoadQueue.scala 163:19:@5607.4]
  assign storeAddrNotKnownFlags_7_5 = _T_5782 & entriesToCheck_7_5; // @[LoadQueue.scala 163:19:@5609.4]
  assign storeAddrNotKnownFlags_7_6 = _T_5785 & entriesToCheck_7_6; // @[LoadQueue.scala 163:19:@5611.4]
  assign storeAddrNotKnownFlags_7_7 = _T_5788 & entriesToCheck_7_7; // @[LoadQueue.scala 163:19:@5613.4]
  assign _T_6122 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0}; // @[Mux.scala 19:72:@5720.4]
  assign _T_6124 = _T_1513 ? _T_6122 : 8'h0; // @[Mux.scala 19:72:@5721.4]
  assign _T_6131 = {conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1}; // @[Mux.scala 19:72:@5728.4]
  assign _T_6133 = _T_1514 ? _T_6131 : 8'h0; // @[Mux.scala 19:72:@5729.4]
  assign _T_6140 = {conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2}; // @[Mux.scala 19:72:@5736.4]
  assign _T_6142 = _T_1515 ? _T_6140 : 8'h0; // @[Mux.scala 19:72:@5737.4]
  assign _T_6149 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3}; // @[Mux.scala 19:72:@5744.4]
  assign _T_6151 = _T_1516 ? _T_6149 : 8'h0; // @[Mux.scala 19:72:@5745.4]
  assign _T_6158 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4}; // @[Mux.scala 19:72:@5752.4]
  assign _T_6160 = _T_1517 ? _T_6158 : 8'h0; // @[Mux.scala 19:72:@5753.4]
  assign _T_6167 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6,conflict_0_5}; // @[Mux.scala 19:72:@5760.4]
  assign _T_6169 = _T_1518 ? _T_6167 : 8'h0; // @[Mux.scala 19:72:@5761.4]
  assign _T_6176 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7,conflict_0_6}; // @[Mux.scala 19:72:@5768.4]
  assign _T_6178 = _T_1519 ? _T_6176 : 8'h0; // @[Mux.scala 19:72:@5769.4]
  assign _T_6185 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_7}; // @[Mux.scala 19:72:@5776.4]
  assign _T_6187 = _T_1520 ? _T_6185 : 8'h0; // @[Mux.scala 19:72:@5777.4]
  assign _T_6188 = _T_6124 | _T_6133; // @[Mux.scala 19:72:@5778.4]
  assign _T_6189 = _T_6188 | _T_6142; // @[Mux.scala 19:72:@5779.4]
  assign _T_6190 = _T_6189 | _T_6151; // @[Mux.scala 19:72:@5780.4]
  assign _T_6191 = _T_6190 | _T_6160; // @[Mux.scala 19:72:@5781.4]
  assign _T_6192 = _T_6191 | _T_6169; // @[Mux.scala 19:72:@5782.4]
  assign _T_6193 = _T_6192 | _T_6178; // @[Mux.scala 19:72:@5783.4]
  assign _T_6194 = _T_6193 | _T_6187; // @[Mux.scala 19:72:@5784.4]
  assign _T_6436 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0}; // @[Mux.scala 19:72:@5902.4]
  assign _T_6438 = _T_1513 ? _T_6436 : 8'h0; // @[Mux.scala 19:72:@5903.4]
  assign _T_6445 = {conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1}; // @[Mux.scala 19:72:@5910.4]
  assign _T_6447 = _T_1514 ? _T_6445 : 8'h0; // @[Mux.scala 19:72:@5911.4]
  assign _T_6454 = {conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2}; // @[Mux.scala 19:72:@5918.4]
  assign _T_6456 = _T_1515 ? _T_6454 : 8'h0; // @[Mux.scala 19:72:@5919.4]
  assign _T_6463 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3}; // @[Mux.scala 19:72:@5926.4]
  assign _T_6465 = _T_1516 ? _T_6463 : 8'h0; // @[Mux.scala 19:72:@5927.4]
  assign _T_6472 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4}; // @[Mux.scala 19:72:@5934.4]
  assign _T_6474 = _T_1517 ? _T_6472 : 8'h0; // @[Mux.scala 19:72:@5935.4]
  assign _T_6481 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6,conflict_1_5}; // @[Mux.scala 19:72:@5942.4]
  assign _T_6483 = _T_1518 ? _T_6481 : 8'h0; // @[Mux.scala 19:72:@5943.4]
  assign _T_6490 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7,conflict_1_6}; // @[Mux.scala 19:72:@5950.4]
  assign _T_6492 = _T_1519 ? _T_6490 : 8'h0; // @[Mux.scala 19:72:@5951.4]
  assign _T_6499 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_7}; // @[Mux.scala 19:72:@5958.4]
  assign _T_6501 = _T_1520 ? _T_6499 : 8'h0; // @[Mux.scala 19:72:@5959.4]
  assign _T_6502 = _T_6438 | _T_6447; // @[Mux.scala 19:72:@5960.4]
  assign _T_6503 = _T_6502 | _T_6456; // @[Mux.scala 19:72:@5961.4]
  assign _T_6504 = _T_6503 | _T_6465; // @[Mux.scala 19:72:@5962.4]
  assign _T_6505 = _T_6504 | _T_6474; // @[Mux.scala 19:72:@5963.4]
  assign _T_6506 = _T_6505 | _T_6483; // @[Mux.scala 19:72:@5964.4]
  assign _T_6507 = _T_6506 | _T_6492; // @[Mux.scala 19:72:@5965.4]
  assign _T_6508 = _T_6507 | _T_6501; // @[Mux.scala 19:72:@5966.4]
  assign _T_6750 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0}; // @[Mux.scala 19:72:@6084.4]
  assign _T_6752 = _T_1513 ? _T_6750 : 8'h0; // @[Mux.scala 19:72:@6085.4]
  assign _T_6759 = {conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1}; // @[Mux.scala 19:72:@6092.4]
  assign _T_6761 = _T_1514 ? _T_6759 : 8'h0; // @[Mux.scala 19:72:@6093.4]
  assign _T_6768 = {conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2}; // @[Mux.scala 19:72:@6100.4]
  assign _T_6770 = _T_1515 ? _T_6768 : 8'h0; // @[Mux.scala 19:72:@6101.4]
  assign _T_6777 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3}; // @[Mux.scala 19:72:@6108.4]
  assign _T_6779 = _T_1516 ? _T_6777 : 8'h0; // @[Mux.scala 19:72:@6109.4]
  assign _T_6786 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4}; // @[Mux.scala 19:72:@6116.4]
  assign _T_6788 = _T_1517 ? _T_6786 : 8'h0; // @[Mux.scala 19:72:@6117.4]
  assign _T_6795 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6,conflict_2_5}; // @[Mux.scala 19:72:@6124.4]
  assign _T_6797 = _T_1518 ? _T_6795 : 8'h0; // @[Mux.scala 19:72:@6125.4]
  assign _T_6804 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7,conflict_2_6}; // @[Mux.scala 19:72:@6132.4]
  assign _T_6806 = _T_1519 ? _T_6804 : 8'h0; // @[Mux.scala 19:72:@6133.4]
  assign _T_6813 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_7}; // @[Mux.scala 19:72:@6140.4]
  assign _T_6815 = _T_1520 ? _T_6813 : 8'h0; // @[Mux.scala 19:72:@6141.4]
  assign _T_6816 = _T_6752 | _T_6761; // @[Mux.scala 19:72:@6142.4]
  assign _T_6817 = _T_6816 | _T_6770; // @[Mux.scala 19:72:@6143.4]
  assign _T_6818 = _T_6817 | _T_6779; // @[Mux.scala 19:72:@6144.4]
  assign _T_6819 = _T_6818 | _T_6788; // @[Mux.scala 19:72:@6145.4]
  assign _T_6820 = _T_6819 | _T_6797; // @[Mux.scala 19:72:@6146.4]
  assign _T_6821 = _T_6820 | _T_6806; // @[Mux.scala 19:72:@6147.4]
  assign _T_6822 = _T_6821 | _T_6815; // @[Mux.scala 19:72:@6148.4]
  assign _T_7064 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0}; // @[Mux.scala 19:72:@6266.4]
  assign _T_7066 = _T_1513 ? _T_7064 : 8'h0; // @[Mux.scala 19:72:@6267.4]
  assign _T_7073 = {conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1}; // @[Mux.scala 19:72:@6274.4]
  assign _T_7075 = _T_1514 ? _T_7073 : 8'h0; // @[Mux.scala 19:72:@6275.4]
  assign _T_7082 = {conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2}; // @[Mux.scala 19:72:@6282.4]
  assign _T_7084 = _T_1515 ? _T_7082 : 8'h0; // @[Mux.scala 19:72:@6283.4]
  assign _T_7091 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3}; // @[Mux.scala 19:72:@6290.4]
  assign _T_7093 = _T_1516 ? _T_7091 : 8'h0; // @[Mux.scala 19:72:@6291.4]
  assign _T_7100 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4}; // @[Mux.scala 19:72:@6298.4]
  assign _T_7102 = _T_1517 ? _T_7100 : 8'h0; // @[Mux.scala 19:72:@6299.4]
  assign _T_7109 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6,conflict_3_5}; // @[Mux.scala 19:72:@6306.4]
  assign _T_7111 = _T_1518 ? _T_7109 : 8'h0; // @[Mux.scala 19:72:@6307.4]
  assign _T_7118 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7,conflict_3_6}; // @[Mux.scala 19:72:@6314.4]
  assign _T_7120 = _T_1519 ? _T_7118 : 8'h0; // @[Mux.scala 19:72:@6315.4]
  assign _T_7127 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_7}; // @[Mux.scala 19:72:@6322.4]
  assign _T_7129 = _T_1520 ? _T_7127 : 8'h0; // @[Mux.scala 19:72:@6323.4]
  assign _T_7130 = _T_7066 | _T_7075; // @[Mux.scala 19:72:@6324.4]
  assign _T_7131 = _T_7130 | _T_7084; // @[Mux.scala 19:72:@6325.4]
  assign _T_7132 = _T_7131 | _T_7093; // @[Mux.scala 19:72:@6326.4]
  assign _T_7133 = _T_7132 | _T_7102; // @[Mux.scala 19:72:@6327.4]
  assign _T_7134 = _T_7133 | _T_7111; // @[Mux.scala 19:72:@6328.4]
  assign _T_7135 = _T_7134 | _T_7120; // @[Mux.scala 19:72:@6329.4]
  assign _T_7136 = _T_7135 | _T_7129; // @[Mux.scala 19:72:@6330.4]
  assign _T_7378 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0}; // @[Mux.scala 19:72:@6448.4]
  assign _T_7380 = _T_1513 ? _T_7378 : 8'h0; // @[Mux.scala 19:72:@6449.4]
  assign _T_7387 = {conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1}; // @[Mux.scala 19:72:@6456.4]
  assign _T_7389 = _T_1514 ? _T_7387 : 8'h0; // @[Mux.scala 19:72:@6457.4]
  assign _T_7396 = {conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2}; // @[Mux.scala 19:72:@6464.4]
  assign _T_7398 = _T_1515 ? _T_7396 : 8'h0; // @[Mux.scala 19:72:@6465.4]
  assign _T_7405 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3}; // @[Mux.scala 19:72:@6472.4]
  assign _T_7407 = _T_1516 ? _T_7405 : 8'h0; // @[Mux.scala 19:72:@6473.4]
  assign _T_7414 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4}; // @[Mux.scala 19:72:@6480.4]
  assign _T_7416 = _T_1517 ? _T_7414 : 8'h0; // @[Mux.scala 19:72:@6481.4]
  assign _T_7423 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6,conflict_4_5}; // @[Mux.scala 19:72:@6488.4]
  assign _T_7425 = _T_1518 ? _T_7423 : 8'h0; // @[Mux.scala 19:72:@6489.4]
  assign _T_7432 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7,conflict_4_6}; // @[Mux.scala 19:72:@6496.4]
  assign _T_7434 = _T_1519 ? _T_7432 : 8'h0; // @[Mux.scala 19:72:@6497.4]
  assign _T_7441 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_7}; // @[Mux.scala 19:72:@6504.4]
  assign _T_7443 = _T_1520 ? _T_7441 : 8'h0; // @[Mux.scala 19:72:@6505.4]
  assign _T_7444 = _T_7380 | _T_7389; // @[Mux.scala 19:72:@6506.4]
  assign _T_7445 = _T_7444 | _T_7398; // @[Mux.scala 19:72:@6507.4]
  assign _T_7446 = _T_7445 | _T_7407; // @[Mux.scala 19:72:@6508.4]
  assign _T_7447 = _T_7446 | _T_7416; // @[Mux.scala 19:72:@6509.4]
  assign _T_7448 = _T_7447 | _T_7425; // @[Mux.scala 19:72:@6510.4]
  assign _T_7449 = _T_7448 | _T_7434; // @[Mux.scala 19:72:@6511.4]
  assign _T_7450 = _T_7449 | _T_7443; // @[Mux.scala 19:72:@6512.4]
  assign _T_7692 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0}; // @[Mux.scala 19:72:@6630.4]
  assign _T_7694 = _T_1513 ? _T_7692 : 8'h0; // @[Mux.scala 19:72:@6631.4]
  assign _T_7701 = {conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1}; // @[Mux.scala 19:72:@6638.4]
  assign _T_7703 = _T_1514 ? _T_7701 : 8'h0; // @[Mux.scala 19:72:@6639.4]
  assign _T_7710 = {conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2}; // @[Mux.scala 19:72:@6646.4]
  assign _T_7712 = _T_1515 ? _T_7710 : 8'h0; // @[Mux.scala 19:72:@6647.4]
  assign _T_7719 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3}; // @[Mux.scala 19:72:@6654.4]
  assign _T_7721 = _T_1516 ? _T_7719 : 8'h0; // @[Mux.scala 19:72:@6655.4]
  assign _T_7728 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4}; // @[Mux.scala 19:72:@6662.4]
  assign _T_7730 = _T_1517 ? _T_7728 : 8'h0; // @[Mux.scala 19:72:@6663.4]
  assign _T_7737 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6,conflict_5_5}; // @[Mux.scala 19:72:@6670.4]
  assign _T_7739 = _T_1518 ? _T_7737 : 8'h0; // @[Mux.scala 19:72:@6671.4]
  assign _T_7746 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7,conflict_5_6}; // @[Mux.scala 19:72:@6678.4]
  assign _T_7748 = _T_1519 ? _T_7746 : 8'h0; // @[Mux.scala 19:72:@6679.4]
  assign _T_7755 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_7}; // @[Mux.scala 19:72:@6686.4]
  assign _T_7757 = _T_1520 ? _T_7755 : 8'h0; // @[Mux.scala 19:72:@6687.4]
  assign _T_7758 = _T_7694 | _T_7703; // @[Mux.scala 19:72:@6688.4]
  assign _T_7759 = _T_7758 | _T_7712; // @[Mux.scala 19:72:@6689.4]
  assign _T_7760 = _T_7759 | _T_7721; // @[Mux.scala 19:72:@6690.4]
  assign _T_7761 = _T_7760 | _T_7730; // @[Mux.scala 19:72:@6691.4]
  assign _T_7762 = _T_7761 | _T_7739; // @[Mux.scala 19:72:@6692.4]
  assign _T_7763 = _T_7762 | _T_7748; // @[Mux.scala 19:72:@6693.4]
  assign _T_7764 = _T_7763 | _T_7757; // @[Mux.scala 19:72:@6694.4]
  assign _T_8006 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0}; // @[Mux.scala 19:72:@6812.4]
  assign _T_8008 = _T_1513 ? _T_8006 : 8'h0; // @[Mux.scala 19:72:@6813.4]
  assign _T_8015 = {conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1}; // @[Mux.scala 19:72:@6820.4]
  assign _T_8017 = _T_1514 ? _T_8015 : 8'h0; // @[Mux.scala 19:72:@6821.4]
  assign _T_8024 = {conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2}; // @[Mux.scala 19:72:@6828.4]
  assign _T_8026 = _T_1515 ? _T_8024 : 8'h0; // @[Mux.scala 19:72:@6829.4]
  assign _T_8033 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3}; // @[Mux.scala 19:72:@6836.4]
  assign _T_8035 = _T_1516 ? _T_8033 : 8'h0; // @[Mux.scala 19:72:@6837.4]
  assign _T_8042 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4}; // @[Mux.scala 19:72:@6844.4]
  assign _T_8044 = _T_1517 ? _T_8042 : 8'h0; // @[Mux.scala 19:72:@6845.4]
  assign _T_8051 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6,conflict_6_5}; // @[Mux.scala 19:72:@6852.4]
  assign _T_8053 = _T_1518 ? _T_8051 : 8'h0; // @[Mux.scala 19:72:@6853.4]
  assign _T_8060 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7,conflict_6_6}; // @[Mux.scala 19:72:@6860.4]
  assign _T_8062 = _T_1519 ? _T_8060 : 8'h0; // @[Mux.scala 19:72:@6861.4]
  assign _T_8069 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_7}; // @[Mux.scala 19:72:@6868.4]
  assign _T_8071 = _T_1520 ? _T_8069 : 8'h0; // @[Mux.scala 19:72:@6869.4]
  assign _T_8072 = _T_8008 | _T_8017; // @[Mux.scala 19:72:@6870.4]
  assign _T_8073 = _T_8072 | _T_8026; // @[Mux.scala 19:72:@6871.4]
  assign _T_8074 = _T_8073 | _T_8035; // @[Mux.scala 19:72:@6872.4]
  assign _T_8075 = _T_8074 | _T_8044; // @[Mux.scala 19:72:@6873.4]
  assign _T_8076 = _T_8075 | _T_8053; // @[Mux.scala 19:72:@6874.4]
  assign _T_8077 = _T_8076 | _T_8062; // @[Mux.scala 19:72:@6875.4]
  assign _T_8078 = _T_8077 | _T_8071; // @[Mux.scala 19:72:@6876.4]
  assign _T_8320 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0}; // @[Mux.scala 19:72:@6994.4]
  assign _T_8322 = _T_1513 ? _T_8320 : 8'h0; // @[Mux.scala 19:72:@6995.4]
  assign _T_8329 = {conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1}; // @[Mux.scala 19:72:@7002.4]
  assign _T_8331 = _T_1514 ? _T_8329 : 8'h0; // @[Mux.scala 19:72:@7003.4]
  assign _T_8338 = {conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2}; // @[Mux.scala 19:72:@7010.4]
  assign _T_8340 = _T_1515 ? _T_8338 : 8'h0; // @[Mux.scala 19:72:@7011.4]
  assign _T_8347 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3}; // @[Mux.scala 19:72:@7018.4]
  assign _T_8349 = _T_1516 ? _T_8347 : 8'h0; // @[Mux.scala 19:72:@7019.4]
  assign _T_8356 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4}; // @[Mux.scala 19:72:@7026.4]
  assign _T_8358 = _T_1517 ? _T_8356 : 8'h0; // @[Mux.scala 19:72:@7027.4]
  assign _T_8365 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6,conflict_7_5}; // @[Mux.scala 19:72:@7034.4]
  assign _T_8367 = _T_1518 ? _T_8365 : 8'h0; // @[Mux.scala 19:72:@7035.4]
  assign _T_8374 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7,conflict_7_6}; // @[Mux.scala 19:72:@7042.4]
  assign _T_8376 = _T_1519 ? _T_8374 : 8'h0; // @[Mux.scala 19:72:@7043.4]
  assign _T_8383 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_7}; // @[Mux.scala 19:72:@7050.4]
  assign _T_8385 = _T_1520 ? _T_8383 : 8'h0; // @[Mux.scala 19:72:@7051.4]
  assign _T_8386 = _T_8322 | _T_8331; // @[Mux.scala 19:72:@7052.4]
  assign _T_8387 = _T_8386 | _T_8340; // @[Mux.scala 19:72:@7053.4]
  assign _T_8388 = _T_8387 | _T_8349; // @[Mux.scala 19:72:@7054.4]
  assign _T_8389 = _T_8388 | _T_8358; // @[Mux.scala 19:72:@7055.4]
  assign _T_8390 = _T_8389 | _T_8367; // @[Mux.scala 19:72:@7056.4]
  assign _T_8391 = _T_8390 | _T_8376; // @[Mux.scala 19:72:@7057.4]
  assign _T_8392 = _T_8391 | _T_8385; // @[Mux.scala 19:72:@7058.4]
  assign _T_14502 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0}; // @[Mux.scala 19:72:@7306.4]
  assign _T_14504 = _T_1513 ? _T_14502 : 8'h0; // @[Mux.scala 19:72:@7307.4]
  assign _T_14511 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1}; // @[Mux.scala 19:72:@7314.4]
  assign _T_14513 = _T_1514 ? _T_14511 : 8'h0; // @[Mux.scala 19:72:@7315.4]
  assign _T_14520 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2}; // @[Mux.scala 19:72:@7322.4]
  assign _T_14522 = _T_1515 ? _T_14520 : 8'h0; // @[Mux.scala 19:72:@7323.4]
  assign _T_14529 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3}; // @[Mux.scala 19:72:@7330.4]
  assign _T_14531 = _T_1516 ? _T_14529 : 8'h0; // @[Mux.scala 19:72:@7331.4]
  assign _T_14538 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4}; // @[Mux.scala 19:72:@7338.4]
  assign _T_14540 = _T_1517 ? _T_14538 : 8'h0; // @[Mux.scala 19:72:@7339.4]
  assign _T_14547 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5}; // @[Mux.scala 19:72:@7346.4]
  assign _T_14549 = _T_1518 ? _T_14547 : 8'h0; // @[Mux.scala 19:72:@7347.4]
  assign _T_14556 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6}; // @[Mux.scala 19:72:@7354.4]
  assign _T_14558 = _T_1519 ? _T_14556 : 8'h0; // @[Mux.scala 19:72:@7355.4]
  assign _T_14565 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_7}; // @[Mux.scala 19:72:@7362.4]
  assign _T_14567 = _T_1520 ? _T_14565 : 8'h0; // @[Mux.scala 19:72:@7363.4]
  assign _T_14568 = _T_14504 | _T_14513; // @[Mux.scala 19:72:@7364.4]
  assign _T_14569 = _T_14568 | _T_14522; // @[Mux.scala 19:72:@7365.4]
  assign _T_14570 = _T_14569 | _T_14531; // @[Mux.scala 19:72:@7366.4]
  assign _T_14571 = _T_14570 | _T_14540; // @[Mux.scala 19:72:@7367.4]
  assign _T_14572 = _T_14571 | _T_14549; // @[Mux.scala 19:72:@7368.4]
  assign _T_14573 = _T_14572 | _T_14558; // @[Mux.scala 19:72:@7369.4]
  assign _T_14574 = _T_14573 | _T_14567; // @[Mux.scala 19:72:@7370.4]
  assign _T_14816 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0}; // @[Mux.scala 19:72:@7488.4]
  assign _T_14818 = _T_1513 ? _T_14816 : 8'h0; // @[Mux.scala 19:72:@7489.4]
  assign _T_14825 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1}; // @[Mux.scala 19:72:@7496.4]
  assign _T_14827 = _T_1514 ? _T_14825 : 8'h0; // @[Mux.scala 19:72:@7497.4]
  assign _T_14834 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2}; // @[Mux.scala 19:72:@7504.4]
  assign _T_14836 = _T_1515 ? _T_14834 : 8'h0; // @[Mux.scala 19:72:@7505.4]
  assign _T_14843 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3}; // @[Mux.scala 19:72:@7512.4]
  assign _T_14845 = _T_1516 ? _T_14843 : 8'h0; // @[Mux.scala 19:72:@7513.4]
  assign _T_14852 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4}; // @[Mux.scala 19:72:@7520.4]
  assign _T_14854 = _T_1517 ? _T_14852 : 8'h0; // @[Mux.scala 19:72:@7521.4]
  assign _T_14861 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5}; // @[Mux.scala 19:72:@7528.4]
  assign _T_14863 = _T_1518 ? _T_14861 : 8'h0; // @[Mux.scala 19:72:@7529.4]
  assign _T_14870 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6}; // @[Mux.scala 19:72:@7536.4]
  assign _T_14872 = _T_1519 ? _T_14870 : 8'h0; // @[Mux.scala 19:72:@7537.4]
  assign _T_14879 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_7}; // @[Mux.scala 19:72:@7544.4]
  assign _T_14881 = _T_1520 ? _T_14879 : 8'h0; // @[Mux.scala 19:72:@7545.4]
  assign _T_14882 = _T_14818 | _T_14827; // @[Mux.scala 19:72:@7546.4]
  assign _T_14883 = _T_14882 | _T_14836; // @[Mux.scala 19:72:@7547.4]
  assign _T_14884 = _T_14883 | _T_14845; // @[Mux.scala 19:72:@7548.4]
  assign _T_14885 = _T_14884 | _T_14854; // @[Mux.scala 19:72:@7549.4]
  assign _T_14886 = _T_14885 | _T_14863; // @[Mux.scala 19:72:@7550.4]
  assign _T_14887 = _T_14886 | _T_14872; // @[Mux.scala 19:72:@7551.4]
  assign _T_14888 = _T_14887 | _T_14881; // @[Mux.scala 19:72:@7552.4]
  assign _T_15130 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0}; // @[Mux.scala 19:72:@7670.4]
  assign _T_15132 = _T_1513 ? _T_15130 : 8'h0; // @[Mux.scala 19:72:@7671.4]
  assign _T_15139 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1}; // @[Mux.scala 19:72:@7678.4]
  assign _T_15141 = _T_1514 ? _T_15139 : 8'h0; // @[Mux.scala 19:72:@7679.4]
  assign _T_15148 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2}; // @[Mux.scala 19:72:@7686.4]
  assign _T_15150 = _T_1515 ? _T_15148 : 8'h0; // @[Mux.scala 19:72:@7687.4]
  assign _T_15157 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3}; // @[Mux.scala 19:72:@7694.4]
  assign _T_15159 = _T_1516 ? _T_15157 : 8'h0; // @[Mux.scala 19:72:@7695.4]
  assign _T_15166 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4}; // @[Mux.scala 19:72:@7702.4]
  assign _T_15168 = _T_1517 ? _T_15166 : 8'h0; // @[Mux.scala 19:72:@7703.4]
  assign _T_15175 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5}; // @[Mux.scala 19:72:@7710.4]
  assign _T_15177 = _T_1518 ? _T_15175 : 8'h0; // @[Mux.scala 19:72:@7711.4]
  assign _T_15184 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6}; // @[Mux.scala 19:72:@7718.4]
  assign _T_15186 = _T_1519 ? _T_15184 : 8'h0; // @[Mux.scala 19:72:@7719.4]
  assign _T_15193 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_7}; // @[Mux.scala 19:72:@7726.4]
  assign _T_15195 = _T_1520 ? _T_15193 : 8'h0; // @[Mux.scala 19:72:@7727.4]
  assign _T_15196 = _T_15132 | _T_15141; // @[Mux.scala 19:72:@7728.4]
  assign _T_15197 = _T_15196 | _T_15150; // @[Mux.scala 19:72:@7729.4]
  assign _T_15198 = _T_15197 | _T_15159; // @[Mux.scala 19:72:@7730.4]
  assign _T_15199 = _T_15198 | _T_15168; // @[Mux.scala 19:72:@7731.4]
  assign _T_15200 = _T_15199 | _T_15177; // @[Mux.scala 19:72:@7732.4]
  assign _T_15201 = _T_15200 | _T_15186; // @[Mux.scala 19:72:@7733.4]
  assign _T_15202 = _T_15201 | _T_15195; // @[Mux.scala 19:72:@7734.4]
  assign _T_15444 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0}; // @[Mux.scala 19:72:@7852.4]
  assign _T_15446 = _T_1513 ? _T_15444 : 8'h0; // @[Mux.scala 19:72:@7853.4]
  assign _T_15453 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1}; // @[Mux.scala 19:72:@7860.4]
  assign _T_15455 = _T_1514 ? _T_15453 : 8'h0; // @[Mux.scala 19:72:@7861.4]
  assign _T_15462 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2}; // @[Mux.scala 19:72:@7868.4]
  assign _T_15464 = _T_1515 ? _T_15462 : 8'h0; // @[Mux.scala 19:72:@7869.4]
  assign _T_15471 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3}; // @[Mux.scala 19:72:@7876.4]
  assign _T_15473 = _T_1516 ? _T_15471 : 8'h0; // @[Mux.scala 19:72:@7877.4]
  assign _T_15480 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4}; // @[Mux.scala 19:72:@7884.4]
  assign _T_15482 = _T_1517 ? _T_15480 : 8'h0; // @[Mux.scala 19:72:@7885.4]
  assign _T_15489 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5}; // @[Mux.scala 19:72:@7892.4]
  assign _T_15491 = _T_1518 ? _T_15489 : 8'h0; // @[Mux.scala 19:72:@7893.4]
  assign _T_15498 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6}; // @[Mux.scala 19:72:@7900.4]
  assign _T_15500 = _T_1519 ? _T_15498 : 8'h0; // @[Mux.scala 19:72:@7901.4]
  assign _T_15507 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_7}; // @[Mux.scala 19:72:@7908.4]
  assign _T_15509 = _T_1520 ? _T_15507 : 8'h0; // @[Mux.scala 19:72:@7909.4]
  assign _T_15510 = _T_15446 | _T_15455; // @[Mux.scala 19:72:@7910.4]
  assign _T_15511 = _T_15510 | _T_15464; // @[Mux.scala 19:72:@7911.4]
  assign _T_15512 = _T_15511 | _T_15473; // @[Mux.scala 19:72:@7912.4]
  assign _T_15513 = _T_15512 | _T_15482; // @[Mux.scala 19:72:@7913.4]
  assign _T_15514 = _T_15513 | _T_15491; // @[Mux.scala 19:72:@7914.4]
  assign _T_15515 = _T_15514 | _T_15500; // @[Mux.scala 19:72:@7915.4]
  assign _T_15516 = _T_15515 | _T_15509; // @[Mux.scala 19:72:@7916.4]
  assign _T_15758 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0}; // @[Mux.scala 19:72:@8034.4]
  assign _T_15760 = _T_1513 ? _T_15758 : 8'h0; // @[Mux.scala 19:72:@8035.4]
  assign _T_15767 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1}; // @[Mux.scala 19:72:@8042.4]
  assign _T_15769 = _T_1514 ? _T_15767 : 8'h0; // @[Mux.scala 19:72:@8043.4]
  assign _T_15776 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2}; // @[Mux.scala 19:72:@8050.4]
  assign _T_15778 = _T_1515 ? _T_15776 : 8'h0; // @[Mux.scala 19:72:@8051.4]
  assign _T_15785 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3}; // @[Mux.scala 19:72:@8058.4]
  assign _T_15787 = _T_1516 ? _T_15785 : 8'h0; // @[Mux.scala 19:72:@8059.4]
  assign _T_15794 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4}; // @[Mux.scala 19:72:@8066.4]
  assign _T_15796 = _T_1517 ? _T_15794 : 8'h0; // @[Mux.scala 19:72:@8067.4]
  assign _T_15803 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5}; // @[Mux.scala 19:72:@8074.4]
  assign _T_15805 = _T_1518 ? _T_15803 : 8'h0; // @[Mux.scala 19:72:@8075.4]
  assign _T_15812 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6}; // @[Mux.scala 19:72:@8082.4]
  assign _T_15814 = _T_1519 ? _T_15812 : 8'h0; // @[Mux.scala 19:72:@8083.4]
  assign _T_15821 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_7}; // @[Mux.scala 19:72:@8090.4]
  assign _T_15823 = _T_1520 ? _T_15821 : 8'h0; // @[Mux.scala 19:72:@8091.4]
  assign _T_15824 = _T_15760 | _T_15769; // @[Mux.scala 19:72:@8092.4]
  assign _T_15825 = _T_15824 | _T_15778; // @[Mux.scala 19:72:@8093.4]
  assign _T_15826 = _T_15825 | _T_15787; // @[Mux.scala 19:72:@8094.4]
  assign _T_15827 = _T_15826 | _T_15796; // @[Mux.scala 19:72:@8095.4]
  assign _T_15828 = _T_15827 | _T_15805; // @[Mux.scala 19:72:@8096.4]
  assign _T_15829 = _T_15828 | _T_15814; // @[Mux.scala 19:72:@8097.4]
  assign _T_15830 = _T_15829 | _T_15823; // @[Mux.scala 19:72:@8098.4]
  assign _T_16072 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0}; // @[Mux.scala 19:72:@8216.4]
  assign _T_16074 = _T_1513 ? _T_16072 : 8'h0; // @[Mux.scala 19:72:@8217.4]
  assign _T_16081 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1}; // @[Mux.scala 19:72:@8224.4]
  assign _T_16083 = _T_1514 ? _T_16081 : 8'h0; // @[Mux.scala 19:72:@8225.4]
  assign _T_16090 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2}; // @[Mux.scala 19:72:@8232.4]
  assign _T_16092 = _T_1515 ? _T_16090 : 8'h0; // @[Mux.scala 19:72:@8233.4]
  assign _T_16099 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3}; // @[Mux.scala 19:72:@8240.4]
  assign _T_16101 = _T_1516 ? _T_16099 : 8'h0; // @[Mux.scala 19:72:@8241.4]
  assign _T_16108 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4}; // @[Mux.scala 19:72:@8248.4]
  assign _T_16110 = _T_1517 ? _T_16108 : 8'h0; // @[Mux.scala 19:72:@8249.4]
  assign _T_16117 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5}; // @[Mux.scala 19:72:@8256.4]
  assign _T_16119 = _T_1518 ? _T_16117 : 8'h0; // @[Mux.scala 19:72:@8257.4]
  assign _T_16126 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6}; // @[Mux.scala 19:72:@8264.4]
  assign _T_16128 = _T_1519 ? _T_16126 : 8'h0; // @[Mux.scala 19:72:@8265.4]
  assign _T_16135 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_7}; // @[Mux.scala 19:72:@8272.4]
  assign _T_16137 = _T_1520 ? _T_16135 : 8'h0; // @[Mux.scala 19:72:@8273.4]
  assign _T_16138 = _T_16074 | _T_16083; // @[Mux.scala 19:72:@8274.4]
  assign _T_16139 = _T_16138 | _T_16092; // @[Mux.scala 19:72:@8275.4]
  assign _T_16140 = _T_16139 | _T_16101; // @[Mux.scala 19:72:@8276.4]
  assign _T_16141 = _T_16140 | _T_16110; // @[Mux.scala 19:72:@8277.4]
  assign _T_16142 = _T_16141 | _T_16119; // @[Mux.scala 19:72:@8278.4]
  assign _T_16143 = _T_16142 | _T_16128; // @[Mux.scala 19:72:@8279.4]
  assign _T_16144 = _T_16143 | _T_16137; // @[Mux.scala 19:72:@8280.4]
  assign _T_16386 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0}; // @[Mux.scala 19:72:@8398.4]
  assign _T_16388 = _T_1513 ? _T_16386 : 8'h0; // @[Mux.scala 19:72:@8399.4]
  assign _T_16395 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1}; // @[Mux.scala 19:72:@8406.4]
  assign _T_16397 = _T_1514 ? _T_16395 : 8'h0; // @[Mux.scala 19:72:@8407.4]
  assign _T_16404 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2}; // @[Mux.scala 19:72:@8414.4]
  assign _T_16406 = _T_1515 ? _T_16404 : 8'h0; // @[Mux.scala 19:72:@8415.4]
  assign _T_16413 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3}; // @[Mux.scala 19:72:@8422.4]
  assign _T_16415 = _T_1516 ? _T_16413 : 8'h0; // @[Mux.scala 19:72:@8423.4]
  assign _T_16422 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4}; // @[Mux.scala 19:72:@8430.4]
  assign _T_16424 = _T_1517 ? _T_16422 : 8'h0; // @[Mux.scala 19:72:@8431.4]
  assign _T_16431 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5}; // @[Mux.scala 19:72:@8438.4]
  assign _T_16433 = _T_1518 ? _T_16431 : 8'h0; // @[Mux.scala 19:72:@8439.4]
  assign _T_16440 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6}; // @[Mux.scala 19:72:@8446.4]
  assign _T_16442 = _T_1519 ? _T_16440 : 8'h0; // @[Mux.scala 19:72:@8447.4]
  assign _T_16449 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_7}; // @[Mux.scala 19:72:@8454.4]
  assign _T_16451 = _T_1520 ? _T_16449 : 8'h0; // @[Mux.scala 19:72:@8455.4]
  assign _T_16452 = _T_16388 | _T_16397; // @[Mux.scala 19:72:@8456.4]
  assign _T_16453 = _T_16452 | _T_16406; // @[Mux.scala 19:72:@8457.4]
  assign _T_16454 = _T_16453 | _T_16415; // @[Mux.scala 19:72:@8458.4]
  assign _T_16455 = _T_16454 | _T_16424; // @[Mux.scala 19:72:@8459.4]
  assign _T_16456 = _T_16455 | _T_16433; // @[Mux.scala 19:72:@8460.4]
  assign _T_16457 = _T_16456 | _T_16442; // @[Mux.scala 19:72:@8461.4]
  assign _T_16458 = _T_16457 | _T_16451; // @[Mux.scala 19:72:@8462.4]
  assign _T_16700 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0}; // @[Mux.scala 19:72:@8580.4]
  assign _T_16702 = _T_1513 ? _T_16700 : 8'h0; // @[Mux.scala 19:72:@8581.4]
  assign _T_16709 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1}; // @[Mux.scala 19:72:@8588.4]
  assign _T_16711 = _T_1514 ? _T_16709 : 8'h0; // @[Mux.scala 19:72:@8589.4]
  assign _T_16718 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2}; // @[Mux.scala 19:72:@8596.4]
  assign _T_16720 = _T_1515 ? _T_16718 : 8'h0; // @[Mux.scala 19:72:@8597.4]
  assign _T_16727 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3}; // @[Mux.scala 19:72:@8604.4]
  assign _T_16729 = _T_1516 ? _T_16727 : 8'h0; // @[Mux.scala 19:72:@8605.4]
  assign _T_16736 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4}; // @[Mux.scala 19:72:@8612.4]
  assign _T_16738 = _T_1517 ? _T_16736 : 8'h0; // @[Mux.scala 19:72:@8613.4]
  assign _T_16745 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5}; // @[Mux.scala 19:72:@8620.4]
  assign _T_16747 = _T_1518 ? _T_16745 : 8'h0; // @[Mux.scala 19:72:@8621.4]
  assign _T_16754 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6}; // @[Mux.scala 19:72:@8628.4]
  assign _T_16756 = _T_1519 ? _T_16754 : 8'h0; // @[Mux.scala 19:72:@8629.4]
  assign _T_16763 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_7}; // @[Mux.scala 19:72:@8636.4]
  assign _T_16765 = _T_1520 ? _T_16763 : 8'h0; // @[Mux.scala 19:72:@8637.4]
  assign _T_16766 = _T_16702 | _T_16711; // @[Mux.scala 19:72:@8638.4]
  assign _T_16767 = _T_16766 | _T_16720; // @[Mux.scala 19:72:@8639.4]
  assign _T_16768 = _T_16767 | _T_16729; // @[Mux.scala 19:72:@8640.4]
  assign _T_16769 = _T_16768 | _T_16738; // @[Mux.scala 19:72:@8641.4]
  assign _T_16770 = _T_16769 | _T_16747; // @[Mux.scala 19:72:@8642.4]
  assign _T_16771 = _T_16770 | _T_16756; // @[Mux.scala 19:72:@8643.4]
  assign _T_16772 = _T_16771 | _T_16765; // @[Mux.scala 19:72:@8644.4]
  assign _T_23532 = conflictPReg_0_2 ? 2'h2 : {{1'd0}, conflictPReg_0_1}; // @[LoadQueue.scala 191:60:@8861.4]
  assign _T_23533 = conflictPReg_0_3 ? 2'h3 : _T_23532; // @[LoadQueue.scala 191:60:@8862.4]
  assign _T_23534 = conflictPReg_0_4 ? 3'h4 : {{1'd0}, _T_23533}; // @[LoadQueue.scala 191:60:@8863.4]
  assign _T_23535 = conflictPReg_0_5 ? 3'h5 : _T_23534; // @[LoadQueue.scala 191:60:@8864.4]
  assign _T_23536 = conflictPReg_0_6 ? 3'h6 : _T_23535; // @[LoadQueue.scala 191:60:@8865.4]
  assign _T_23537 = conflictPReg_0_7 ? 3'h7 : _T_23536; // @[LoadQueue.scala 191:60:@8866.4]
  assign _T_23540 = conflictPReg_0_0 | conflictPReg_0_1; // @[LoadQueue.scala 192:43:@8868.4]
  assign _T_23541 = _T_23540 | conflictPReg_0_2; // @[LoadQueue.scala 192:43:@8869.4]
  assign _T_23542 = _T_23541 | conflictPReg_0_3; // @[LoadQueue.scala 192:43:@8870.4]
  assign _T_23543 = _T_23542 | conflictPReg_0_4; // @[LoadQueue.scala 192:43:@8871.4]
  assign _T_23544 = _T_23543 | conflictPReg_0_5; // @[LoadQueue.scala 192:43:@8872.4]
  assign _T_23545 = _T_23544 | conflictPReg_0_6; // @[LoadQueue.scala 192:43:@8873.4]
  assign _T_23546 = _T_23545 | conflictPReg_0_7; // @[LoadQueue.scala 192:43:@8874.4]
  assign _GEN_240 = 3'h0 == _T_23537; // @[LoadQueue.scala 193:43:@8876.6]
  assign _GEN_241 = 3'h1 == _T_23537; // @[LoadQueue.scala 193:43:@8876.6]
  assign _GEN_242 = 3'h2 == _T_23537; // @[LoadQueue.scala 193:43:@8876.6]
  assign _GEN_243 = 3'h3 == _T_23537; // @[LoadQueue.scala 193:43:@8876.6]
  assign _GEN_244 = 3'h4 == _T_23537; // @[LoadQueue.scala 193:43:@8876.6]
  assign _GEN_245 = 3'h5 == _T_23537; // @[LoadQueue.scala 193:43:@8876.6]
  assign _GEN_246 = 3'h6 == _T_23537; // @[LoadQueue.scala 193:43:@8876.6]
  assign _GEN_247 = 3'h7 == _T_23537; // @[LoadQueue.scala 193:43:@8876.6]
  assign _GEN_249 = 3'h1 == _T_23537 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8877.6]
  assign _GEN_250 = 3'h2 == _T_23537 ? shiftedStoreDataKnownPReg_2 : _GEN_249; // @[LoadQueue.scala 194:31:@8877.6]
  assign _GEN_251 = 3'h3 == _T_23537 ? shiftedStoreDataKnownPReg_3 : _GEN_250; // @[LoadQueue.scala 194:31:@8877.6]
  assign _GEN_252 = 3'h4 == _T_23537 ? shiftedStoreDataKnownPReg_4 : _GEN_251; // @[LoadQueue.scala 194:31:@8877.6]
  assign _GEN_253 = 3'h5 == _T_23537 ? shiftedStoreDataKnownPReg_5 : _GEN_252; // @[LoadQueue.scala 194:31:@8877.6]
  assign _GEN_254 = 3'h6 == _T_23537 ? shiftedStoreDataKnownPReg_6 : _GEN_253; // @[LoadQueue.scala 194:31:@8877.6]
  assign _GEN_255 = 3'h7 == _T_23537 ? shiftedStoreDataKnownPReg_7 : _GEN_254; // @[LoadQueue.scala 194:31:@8877.6]
  assign _GEN_257 = 3'h1 == _T_23537 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8878.6]
  assign _GEN_258 = 3'h2 == _T_23537 ? shiftedStoreDataQPreg_2 : _GEN_257; // @[LoadQueue.scala 195:31:@8878.6]
  assign _GEN_259 = 3'h3 == _T_23537 ? shiftedStoreDataQPreg_3 : _GEN_258; // @[LoadQueue.scala 195:31:@8878.6]
  assign _GEN_260 = 3'h4 == _T_23537 ? shiftedStoreDataQPreg_4 : _GEN_259; // @[LoadQueue.scala 195:31:@8878.6]
  assign _GEN_261 = 3'h5 == _T_23537 ? shiftedStoreDataQPreg_5 : _GEN_260; // @[LoadQueue.scala 195:31:@8878.6]
  assign _GEN_262 = 3'h6 == _T_23537 ? shiftedStoreDataQPreg_6 : _GEN_261; // @[LoadQueue.scala 195:31:@8878.6]
  assign _GEN_263 = 3'h7 == _T_23537 ? shiftedStoreDataQPreg_7 : _GEN_262; // @[LoadQueue.scala 195:31:@8878.6]
  assign lastConflict_0_0 = _T_23546 ? _GEN_240 : 1'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign lastConflict_0_1 = _T_23546 ? _GEN_241 : 1'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign lastConflict_0_2 = _T_23546 ? _GEN_242 : 1'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign lastConflict_0_3 = _T_23546 ? _GEN_243 : 1'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign lastConflict_0_4 = _T_23546 ? _GEN_244 : 1'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign lastConflict_0_5 = _T_23546 ? _GEN_245 : 1'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign lastConflict_0_6 = _T_23546 ? _GEN_246 : 1'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign lastConflict_0_7 = _T_23546 ? _GEN_247 : 1'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign canBypass_0 = _T_23546 ? _GEN_255 : 1'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign bypassVal_0 = _T_23546 ? _GEN_263 : 32'h0; // @[LoadQueue.scala 192:53:@8875.4]
  assign _T_23612 = conflictPReg_1_2 ? 2'h2 : {{1'd0}, conflictPReg_1_1}; // @[LoadQueue.scala 191:60:@8908.4]
  assign _T_23613 = conflictPReg_1_3 ? 2'h3 : _T_23612; // @[LoadQueue.scala 191:60:@8909.4]
  assign _T_23614 = conflictPReg_1_4 ? 3'h4 : {{1'd0}, _T_23613}; // @[LoadQueue.scala 191:60:@8910.4]
  assign _T_23615 = conflictPReg_1_5 ? 3'h5 : _T_23614; // @[LoadQueue.scala 191:60:@8911.4]
  assign _T_23616 = conflictPReg_1_6 ? 3'h6 : _T_23615; // @[LoadQueue.scala 191:60:@8912.4]
  assign _T_23617 = conflictPReg_1_7 ? 3'h7 : _T_23616; // @[LoadQueue.scala 191:60:@8913.4]
  assign _T_23620 = conflictPReg_1_0 | conflictPReg_1_1; // @[LoadQueue.scala 192:43:@8915.4]
  assign _T_23621 = _T_23620 | conflictPReg_1_2; // @[LoadQueue.scala 192:43:@8916.4]
  assign _T_23622 = _T_23621 | conflictPReg_1_3; // @[LoadQueue.scala 192:43:@8917.4]
  assign _T_23623 = _T_23622 | conflictPReg_1_4; // @[LoadQueue.scala 192:43:@8918.4]
  assign _T_23624 = _T_23623 | conflictPReg_1_5; // @[LoadQueue.scala 192:43:@8919.4]
  assign _T_23625 = _T_23624 | conflictPReg_1_6; // @[LoadQueue.scala 192:43:@8920.4]
  assign _T_23626 = _T_23625 | conflictPReg_1_7; // @[LoadQueue.scala 192:43:@8921.4]
  assign _GEN_274 = 3'h0 == _T_23617; // @[LoadQueue.scala 193:43:@8923.6]
  assign _GEN_275 = 3'h1 == _T_23617; // @[LoadQueue.scala 193:43:@8923.6]
  assign _GEN_276 = 3'h2 == _T_23617; // @[LoadQueue.scala 193:43:@8923.6]
  assign _GEN_277 = 3'h3 == _T_23617; // @[LoadQueue.scala 193:43:@8923.6]
  assign _GEN_278 = 3'h4 == _T_23617; // @[LoadQueue.scala 193:43:@8923.6]
  assign _GEN_279 = 3'h5 == _T_23617; // @[LoadQueue.scala 193:43:@8923.6]
  assign _GEN_280 = 3'h6 == _T_23617; // @[LoadQueue.scala 193:43:@8923.6]
  assign _GEN_281 = 3'h7 == _T_23617; // @[LoadQueue.scala 193:43:@8923.6]
  assign _GEN_283 = 3'h1 == _T_23617 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8924.6]
  assign _GEN_284 = 3'h2 == _T_23617 ? shiftedStoreDataKnownPReg_2 : _GEN_283; // @[LoadQueue.scala 194:31:@8924.6]
  assign _GEN_285 = 3'h3 == _T_23617 ? shiftedStoreDataKnownPReg_3 : _GEN_284; // @[LoadQueue.scala 194:31:@8924.6]
  assign _GEN_286 = 3'h4 == _T_23617 ? shiftedStoreDataKnownPReg_4 : _GEN_285; // @[LoadQueue.scala 194:31:@8924.6]
  assign _GEN_287 = 3'h5 == _T_23617 ? shiftedStoreDataKnownPReg_5 : _GEN_286; // @[LoadQueue.scala 194:31:@8924.6]
  assign _GEN_288 = 3'h6 == _T_23617 ? shiftedStoreDataKnownPReg_6 : _GEN_287; // @[LoadQueue.scala 194:31:@8924.6]
  assign _GEN_289 = 3'h7 == _T_23617 ? shiftedStoreDataKnownPReg_7 : _GEN_288; // @[LoadQueue.scala 194:31:@8924.6]
  assign _GEN_291 = 3'h1 == _T_23617 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8925.6]
  assign _GEN_292 = 3'h2 == _T_23617 ? shiftedStoreDataQPreg_2 : _GEN_291; // @[LoadQueue.scala 195:31:@8925.6]
  assign _GEN_293 = 3'h3 == _T_23617 ? shiftedStoreDataQPreg_3 : _GEN_292; // @[LoadQueue.scala 195:31:@8925.6]
  assign _GEN_294 = 3'h4 == _T_23617 ? shiftedStoreDataQPreg_4 : _GEN_293; // @[LoadQueue.scala 195:31:@8925.6]
  assign _GEN_295 = 3'h5 == _T_23617 ? shiftedStoreDataQPreg_5 : _GEN_294; // @[LoadQueue.scala 195:31:@8925.6]
  assign _GEN_296 = 3'h6 == _T_23617 ? shiftedStoreDataQPreg_6 : _GEN_295; // @[LoadQueue.scala 195:31:@8925.6]
  assign _GEN_297 = 3'h7 == _T_23617 ? shiftedStoreDataQPreg_7 : _GEN_296; // @[LoadQueue.scala 195:31:@8925.6]
  assign lastConflict_1_0 = _T_23626 ? _GEN_274 : 1'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign lastConflict_1_1 = _T_23626 ? _GEN_275 : 1'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign lastConflict_1_2 = _T_23626 ? _GEN_276 : 1'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign lastConflict_1_3 = _T_23626 ? _GEN_277 : 1'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign lastConflict_1_4 = _T_23626 ? _GEN_278 : 1'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign lastConflict_1_5 = _T_23626 ? _GEN_279 : 1'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign lastConflict_1_6 = _T_23626 ? _GEN_280 : 1'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign lastConflict_1_7 = _T_23626 ? _GEN_281 : 1'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign canBypass_1 = _T_23626 ? _GEN_289 : 1'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign bypassVal_1 = _T_23626 ? _GEN_297 : 32'h0; // @[LoadQueue.scala 192:53:@8922.4]
  assign _T_23692 = conflictPReg_2_2 ? 2'h2 : {{1'd0}, conflictPReg_2_1}; // @[LoadQueue.scala 191:60:@8955.4]
  assign _T_23693 = conflictPReg_2_3 ? 2'h3 : _T_23692; // @[LoadQueue.scala 191:60:@8956.4]
  assign _T_23694 = conflictPReg_2_4 ? 3'h4 : {{1'd0}, _T_23693}; // @[LoadQueue.scala 191:60:@8957.4]
  assign _T_23695 = conflictPReg_2_5 ? 3'h5 : _T_23694; // @[LoadQueue.scala 191:60:@8958.4]
  assign _T_23696 = conflictPReg_2_6 ? 3'h6 : _T_23695; // @[LoadQueue.scala 191:60:@8959.4]
  assign _T_23697 = conflictPReg_2_7 ? 3'h7 : _T_23696; // @[LoadQueue.scala 191:60:@8960.4]
  assign _T_23700 = conflictPReg_2_0 | conflictPReg_2_1; // @[LoadQueue.scala 192:43:@8962.4]
  assign _T_23701 = _T_23700 | conflictPReg_2_2; // @[LoadQueue.scala 192:43:@8963.4]
  assign _T_23702 = _T_23701 | conflictPReg_2_3; // @[LoadQueue.scala 192:43:@8964.4]
  assign _T_23703 = _T_23702 | conflictPReg_2_4; // @[LoadQueue.scala 192:43:@8965.4]
  assign _T_23704 = _T_23703 | conflictPReg_2_5; // @[LoadQueue.scala 192:43:@8966.4]
  assign _T_23705 = _T_23704 | conflictPReg_2_6; // @[LoadQueue.scala 192:43:@8967.4]
  assign _T_23706 = _T_23705 | conflictPReg_2_7; // @[LoadQueue.scala 192:43:@8968.4]
  assign _GEN_308 = 3'h0 == _T_23697; // @[LoadQueue.scala 193:43:@8970.6]
  assign _GEN_309 = 3'h1 == _T_23697; // @[LoadQueue.scala 193:43:@8970.6]
  assign _GEN_310 = 3'h2 == _T_23697; // @[LoadQueue.scala 193:43:@8970.6]
  assign _GEN_311 = 3'h3 == _T_23697; // @[LoadQueue.scala 193:43:@8970.6]
  assign _GEN_312 = 3'h4 == _T_23697; // @[LoadQueue.scala 193:43:@8970.6]
  assign _GEN_313 = 3'h5 == _T_23697; // @[LoadQueue.scala 193:43:@8970.6]
  assign _GEN_314 = 3'h6 == _T_23697; // @[LoadQueue.scala 193:43:@8970.6]
  assign _GEN_315 = 3'h7 == _T_23697; // @[LoadQueue.scala 193:43:@8970.6]
  assign _GEN_317 = 3'h1 == _T_23697 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@8971.6]
  assign _GEN_318 = 3'h2 == _T_23697 ? shiftedStoreDataKnownPReg_2 : _GEN_317; // @[LoadQueue.scala 194:31:@8971.6]
  assign _GEN_319 = 3'h3 == _T_23697 ? shiftedStoreDataKnownPReg_3 : _GEN_318; // @[LoadQueue.scala 194:31:@8971.6]
  assign _GEN_320 = 3'h4 == _T_23697 ? shiftedStoreDataKnownPReg_4 : _GEN_319; // @[LoadQueue.scala 194:31:@8971.6]
  assign _GEN_321 = 3'h5 == _T_23697 ? shiftedStoreDataKnownPReg_5 : _GEN_320; // @[LoadQueue.scala 194:31:@8971.6]
  assign _GEN_322 = 3'h6 == _T_23697 ? shiftedStoreDataKnownPReg_6 : _GEN_321; // @[LoadQueue.scala 194:31:@8971.6]
  assign _GEN_323 = 3'h7 == _T_23697 ? shiftedStoreDataKnownPReg_7 : _GEN_322; // @[LoadQueue.scala 194:31:@8971.6]
  assign _GEN_325 = 3'h1 == _T_23697 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@8972.6]
  assign _GEN_326 = 3'h2 == _T_23697 ? shiftedStoreDataQPreg_2 : _GEN_325; // @[LoadQueue.scala 195:31:@8972.6]
  assign _GEN_327 = 3'h3 == _T_23697 ? shiftedStoreDataQPreg_3 : _GEN_326; // @[LoadQueue.scala 195:31:@8972.6]
  assign _GEN_328 = 3'h4 == _T_23697 ? shiftedStoreDataQPreg_4 : _GEN_327; // @[LoadQueue.scala 195:31:@8972.6]
  assign _GEN_329 = 3'h5 == _T_23697 ? shiftedStoreDataQPreg_5 : _GEN_328; // @[LoadQueue.scala 195:31:@8972.6]
  assign _GEN_330 = 3'h6 == _T_23697 ? shiftedStoreDataQPreg_6 : _GEN_329; // @[LoadQueue.scala 195:31:@8972.6]
  assign _GEN_331 = 3'h7 == _T_23697 ? shiftedStoreDataQPreg_7 : _GEN_330; // @[LoadQueue.scala 195:31:@8972.6]
  assign lastConflict_2_0 = _T_23706 ? _GEN_308 : 1'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign lastConflict_2_1 = _T_23706 ? _GEN_309 : 1'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign lastConflict_2_2 = _T_23706 ? _GEN_310 : 1'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign lastConflict_2_3 = _T_23706 ? _GEN_311 : 1'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign lastConflict_2_4 = _T_23706 ? _GEN_312 : 1'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign lastConflict_2_5 = _T_23706 ? _GEN_313 : 1'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign lastConflict_2_6 = _T_23706 ? _GEN_314 : 1'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign lastConflict_2_7 = _T_23706 ? _GEN_315 : 1'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign canBypass_2 = _T_23706 ? _GEN_323 : 1'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign bypassVal_2 = _T_23706 ? _GEN_331 : 32'h0; // @[LoadQueue.scala 192:53:@8969.4]
  assign _T_23772 = conflictPReg_3_2 ? 2'h2 : {{1'd0}, conflictPReg_3_1}; // @[LoadQueue.scala 191:60:@9002.4]
  assign _T_23773 = conflictPReg_3_3 ? 2'h3 : _T_23772; // @[LoadQueue.scala 191:60:@9003.4]
  assign _T_23774 = conflictPReg_3_4 ? 3'h4 : {{1'd0}, _T_23773}; // @[LoadQueue.scala 191:60:@9004.4]
  assign _T_23775 = conflictPReg_3_5 ? 3'h5 : _T_23774; // @[LoadQueue.scala 191:60:@9005.4]
  assign _T_23776 = conflictPReg_3_6 ? 3'h6 : _T_23775; // @[LoadQueue.scala 191:60:@9006.4]
  assign _T_23777 = conflictPReg_3_7 ? 3'h7 : _T_23776; // @[LoadQueue.scala 191:60:@9007.4]
  assign _T_23780 = conflictPReg_3_0 | conflictPReg_3_1; // @[LoadQueue.scala 192:43:@9009.4]
  assign _T_23781 = _T_23780 | conflictPReg_3_2; // @[LoadQueue.scala 192:43:@9010.4]
  assign _T_23782 = _T_23781 | conflictPReg_3_3; // @[LoadQueue.scala 192:43:@9011.4]
  assign _T_23783 = _T_23782 | conflictPReg_3_4; // @[LoadQueue.scala 192:43:@9012.4]
  assign _T_23784 = _T_23783 | conflictPReg_3_5; // @[LoadQueue.scala 192:43:@9013.4]
  assign _T_23785 = _T_23784 | conflictPReg_3_6; // @[LoadQueue.scala 192:43:@9014.4]
  assign _T_23786 = _T_23785 | conflictPReg_3_7; // @[LoadQueue.scala 192:43:@9015.4]
  assign _GEN_342 = 3'h0 == _T_23777; // @[LoadQueue.scala 193:43:@9017.6]
  assign _GEN_343 = 3'h1 == _T_23777; // @[LoadQueue.scala 193:43:@9017.6]
  assign _GEN_344 = 3'h2 == _T_23777; // @[LoadQueue.scala 193:43:@9017.6]
  assign _GEN_345 = 3'h3 == _T_23777; // @[LoadQueue.scala 193:43:@9017.6]
  assign _GEN_346 = 3'h4 == _T_23777; // @[LoadQueue.scala 193:43:@9017.6]
  assign _GEN_347 = 3'h5 == _T_23777; // @[LoadQueue.scala 193:43:@9017.6]
  assign _GEN_348 = 3'h6 == _T_23777; // @[LoadQueue.scala 193:43:@9017.6]
  assign _GEN_349 = 3'h7 == _T_23777; // @[LoadQueue.scala 193:43:@9017.6]
  assign _GEN_351 = 3'h1 == _T_23777 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@9018.6]
  assign _GEN_352 = 3'h2 == _T_23777 ? shiftedStoreDataKnownPReg_2 : _GEN_351; // @[LoadQueue.scala 194:31:@9018.6]
  assign _GEN_353 = 3'h3 == _T_23777 ? shiftedStoreDataKnownPReg_3 : _GEN_352; // @[LoadQueue.scala 194:31:@9018.6]
  assign _GEN_354 = 3'h4 == _T_23777 ? shiftedStoreDataKnownPReg_4 : _GEN_353; // @[LoadQueue.scala 194:31:@9018.6]
  assign _GEN_355 = 3'h5 == _T_23777 ? shiftedStoreDataKnownPReg_5 : _GEN_354; // @[LoadQueue.scala 194:31:@9018.6]
  assign _GEN_356 = 3'h6 == _T_23777 ? shiftedStoreDataKnownPReg_6 : _GEN_355; // @[LoadQueue.scala 194:31:@9018.6]
  assign _GEN_357 = 3'h7 == _T_23777 ? shiftedStoreDataKnownPReg_7 : _GEN_356; // @[LoadQueue.scala 194:31:@9018.6]
  assign _GEN_359 = 3'h1 == _T_23777 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@9019.6]
  assign _GEN_360 = 3'h2 == _T_23777 ? shiftedStoreDataQPreg_2 : _GEN_359; // @[LoadQueue.scala 195:31:@9019.6]
  assign _GEN_361 = 3'h3 == _T_23777 ? shiftedStoreDataQPreg_3 : _GEN_360; // @[LoadQueue.scala 195:31:@9019.6]
  assign _GEN_362 = 3'h4 == _T_23777 ? shiftedStoreDataQPreg_4 : _GEN_361; // @[LoadQueue.scala 195:31:@9019.6]
  assign _GEN_363 = 3'h5 == _T_23777 ? shiftedStoreDataQPreg_5 : _GEN_362; // @[LoadQueue.scala 195:31:@9019.6]
  assign _GEN_364 = 3'h6 == _T_23777 ? shiftedStoreDataQPreg_6 : _GEN_363; // @[LoadQueue.scala 195:31:@9019.6]
  assign _GEN_365 = 3'h7 == _T_23777 ? shiftedStoreDataQPreg_7 : _GEN_364; // @[LoadQueue.scala 195:31:@9019.6]
  assign lastConflict_3_0 = _T_23786 ? _GEN_342 : 1'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign lastConflict_3_1 = _T_23786 ? _GEN_343 : 1'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign lastConflict_3_2 = _T_23786 ? _GEN_344 : 1'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign lastConflict_3_3 = _T_23786 ? _GEN_345 : 1'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign lastConflict_3_4 = _T_23786 ? _GEN_346 : 1'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign lastConflict_3_5 = _T_23786 ? _GEN_347 : 1'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign lastConflict_3_6 = _T_23786 ? _GEN_348 : 1'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign lastConflict_3_7 = _T_23786 ? _GEN_349 : 1'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign canBypass_3 = _T_23786 ? _GEN_357 : 1'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign bypassVal_3 = _T_23786 ? _GEN_365 : 32'h0; // @[LoadQueue.scala 192:53:@9016.4]
  assign _T_23852 = conflictPReg_4_2 ? 2'h2 : {{1'd0}, conflictPReg_4_1}; // @[LoadQueue.scala 191:60:@9049.4]
  assign _T_23853 = conflictPReg_4_3 ? 2'h3 : _T_23852; // @[LoadQueue.scala 191:60:@9050.4]
  assign _T_23854 = conflictPReg_4_4 ? 3'h4 : {{1'd0}, _T_23853}; // @[LoadQueue.scala 191:60:@9051.4]
  assign _T_23855 = conflictPReg_4_5 ? 3'h5 : _T_23854; // @[LoadQueue.scala 191:60:@9052.4]
  assign _T_23856 = conflictPReg_4_6 ? 3'h6 : _T_23855; // @[LoadQueue.scala 191:60:@9053.4]
  assign _T_23857 = conflictPReg_4_7 ? 3'h7 : _T_23856; // @[LoadQueue.scala 191:60:@9054.4]
  assign _T_23860 = conflictPReg_4_0 | conflictPReg_4_1; // @[LoadQueue.scala 192:43:@9056.4]
  assign _T_23861 = _T_23860 | conflictPReg_4_2; // @[LoadQueue.scala 192:43:@9057.4]
  assign _T_23862 = _T_23861 | conflictPReg_4_3; // @[LoadQueue.scala 192:43:@9058.4]
  assign _T_23863 = _T_23862 | conflictPReg_4_4; // @[LoadQueue.scala 192:43:@9059.4]
  assign _T_23864 = _T_23863 | conflictPReg_4_5; // @[LoadQueue.scala 192:43:@9060.4]
  assign _T_23865 = _T_23864 | conflictPReg_4_6; // @[LoadQueue.scala 192:43:@9061.4]
  assign _T_23866 = _T_23865 | conflictPReg_4_7; // @[LoadQueue.scala 192:43:@9062.4]
  assign _GEN_376 = 3'h0 == _T_23857; // @[LoadQueue.scala 193:43:@9064.6]
  assign _GEN_377 = 3'h1 == _T_23857; // @[LoadQueue.scala 193:43:@9064.6]
  assign _GEN_378 = 3'h2 == _T_23857; // @[LoadQueue.scala 193:43:@9064.6]
  assign _GEN_379 = 3'h3 == _T_23857; // @[LoadQueue.scala 193:43:@9064.6]
  assign _GEN_380 = 3'h4 == _T_23857; // @[LoadQueue.scala 193:43:@9064.6]
  assign _GEN_381 = 3'h5 == _T_23857; // @[LoadQueue.scala 193:43:@9064.6]
  assign _GEN_382 = 3'h6 == _T_23857; // @[LoadQueue.scala 193:43:@9064.6]
  assign _GEN_383 = 3'h7 == _T_23857; // @[LoadQueue.scala 193:43:@9064.6]
  assign _GEN_385 = 3'h1 == _T_23857 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@9065.6]
  assign _GEN_386 = 3'h2 == _T_23857 ? shiftedStoreDataKnownPReg_2 : _GEN_385; // @[LoadQueue.scala 194:31:@9065.6]
  assign _GEN_387 = 3'h3 == _T_23857 ? shiftedStoreDataKnownPReg_3 : _GEN_386; // @[LoadQueue.scala 194:31:@9065.6]
  assign _GEN_388 = 3'h4 == _T_23857 ? shiftedStoreDataKnownPReg_4 : _GEN_387; // @[LoadQueue.scala 194:31:@9065.6]
  assign _GEN_389 = 3'h5 == _T_23857 ? shiftedStoreDataKnownPReg_5 : _GEN_388; // @[LoadQueue.scala 194:31:@9065.6]
  assign _GEN_390 = 3'h6 == _T_23857 ? shiftedStoreDataKnownPReg_6 : _GEN_389; // @[LoadQueue.scala 194:31:@9065.6]
  assign _GEN_391 = 3'h7 == _T_23857 ? shiftedStoreDataKnownPReg_7 : _GEN_390; // @[LoadQueue.scala 194:31:@9065.6]
  assign _GEN_393 = 3'h1 == _T_23857 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@9066.6]
  assign _GEN_394 = 3'h2 == _T_23857 ? shiftedStoreDataQPreg_2 : _GEN_393; // @[LoadQueue.scala 195:31:@9066.6]
  assign _GEN_395 = 3'h3 == _T_23857 ? shiftedStoreDataQPreg_3 : _GEN_394; // @[LoadQueue.scala 195:31:@9066.6]
  assign _GEN_396 = 3'h4 == _T_23857 ? shiftedStoreDataQPreg_4 : _GEN_395; // @[LoadQueue.scala 195:31:@9066.6]
  assign _GEN_397 = 3'h5 == _T_23857 ? shiftedStoreDataQPreg_5 : _GEN_396; // @[LoadQueue.scala 195:31:@9066.6]
  assign _GEN_398 = 3'h6 == _T_23857 ? shiftedStoreDataQPreg_6 : _GEN_397; // @[LoadQueue.scala 195:31:@9066.6]
  assign _GEN_399 = 3'h7 == _T_23857 ? shiftedStoreDataQPreg_7 : _GEN_398; // @[LoadQueue.scala 195:31:@9066.6]
  assign lastConflict_4_0 = _T_23866 ? _GEN_376 : 1'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign lastConflict_4_1 = _T_23866 ? _GEN_377 : 1'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign lastConflict_4_2 = _T_23866 ? _GEN_378 : 1'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign lastConflict_4_3 = _T_23866 ? _GEN_379 : 1'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign lastConflict_4_4 = _T_23866 ? _GEN_380 : 1'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign lastConflict_4_5 = _T_23866 ? _GEN_381 : 1'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign lastConflict_4_6 = _T_23866 ? _GEN_382 : 1'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign lastConflict_4_7 = _T_23866 ? _GEN_383 : 1'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign canBypass_4 = _T_23866 ? _GEN_391 : 1'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign bypassVal_4 = _T_23866 ? _GEN_399 : 32'h0; // @[LoadQueue.scala 192:53:@9063.4]
  assign _T_23932 = conflictPReg_5_2 ? 2'h2 : {{1'd0}, conflictPReg_5_1}; // @[LoadQueue.scala 191:60:@9096.4]
  assign _T_23933 = conflictPReg_5_3 ? 2'h3 : _T_23932; // @[LoadQueue.scala 191:60:@9097.4]
  assign _T_23934 = conflictPReg_5_4 ? 3'h4 : {{1'd0}, _T_23933}; // @[LoadQueue.scala 191:60:@9098.4]
  assign _T_23935 = conflictPReg_5_5 ? 3'h5 : _T_23934; // @[LoadQueue.scala 191:60:@9099.4]
  assign _T_23936 = conflictPReg_5_6 ? 3'h6 : _T_23935; // @[LoadQueue.scala 191:60:@9100.4]
  assign _T_23937 = conflictPReg_5_7 ? 3'h7 : _T_23936; // @[LoadQueue.scala 191:60:@9101.4]
  assign _T_23940 = conflictPReg_5_0 | conflictPReg_5_1; // @[LoadQueue.scala 192:43:@9103.4]
  assign _T_23941 = _T_23940 | conflictPReg_5_2; // @[LoadQueue.scala 192:43:@9104.4]
  assign _T_23942 = _T_23941 | conflictPReg_5_3; // @[LoadQueue.scala 192:43:@9105.4]
  assign _T_23943 = _T_23942 | conflictPReg_5_4; // @[LoadQueue.scala 192:43:@9106.4]
  assign _T_23944 = _T_23943 | conflictPReg_5_5; // @[LoadQueue.scala 192:43:@9107.4]
  assign _T_23945 = _T_23944 | conflictPReg_5_6; // @[LoadQueue.scala 192:43:@9108.4]
  assign _T_23946 = _T_23945 | conflictPReg_5_7; // @[LoadQueue.scala 192:43:@9109.4]
  assign _GEN_410 = 3'h0 == _T_23937; // @[LoadQueue.scala 193:43:@9111.6]
  assign _GEN_411 = 3'h1 == _T_23937; // @[LoadQueue.scala 193:43:@9111.6]
  assign _GEN_412 = 3'h2 == _T_23937; // @[LoadQueue.scala 193:43:@9111.6]
  assign _GEN_413 = 3'h3 == _T_23937; // @[LoadQueue.scala 193:43:@9111.6]
  assign _GEN_414 = 3'h4 == _T_23937; // @[LoadQueue.scala 193:43:@9111.6]
  assign _GEN_415 = 3'h5 == _T_23937; // @[LoadQueue.scala 193:43:@9111.6]
  assign _GEN_416 = 3'h6 == _T_23937; // @[LoadQueue.scala 193:43:@9111.6]
  assign _GEN_417 = 3'h7 == _T_23937; // @[LoadQueue.scala 193:43:@9111.6]
  assign _GEN_419 = 3'h1 == _T_23937 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@9112.6]
  assign _GEN_420 = 3'h2 == _T_23937 ? shiftedStoreDataKnownPReg_2 : _GEN_419; // @[LoadQueue.scala 194:31:@9112.6]
  assign _GEN_421 = 3'h3 == _T_23937 ? shiftedStoreDataKnownPReg_3 : _GEN_420; // @[LoadQueue.scala 194:31:@9112.6]
  assign _GEN_422 = 3'h4 == _T_23937 ? shiftedStoreDataKnownPReg_4 : _GEN_421; // @[LoadQueue.scala 194:31:@9112.6]
  assign _GEN_423 = 3'h5 == _T_23937 ? shiftedStoreDataKnownPReg_5 : _GEN_422; // @[LoadQueue.scala 194:31:@9112.6]
  assign _GEN_424 = 3'h6 == _T_23937 ? shiftedStoreDataKnownPReg_6 : _GEN_423; // @[LoadQueue.scala 194:31:@9112.6]
  assign _GEN_425 = 3'h7 == _T_23937 ? shiftedStoreDataKnownPReg_7 : _GEN_424; // @[LoadQueue.scala 194:31:@9112.6]
  assign _GEN_427 = 3'h1 == _T_23937 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@9113.6]
  assign _GEN_428 = 3'h2 == _T_23937 ? shiftedStoreDataQPreg_2 : _GEN_427; // @[LoadQueue.scala 195:31:@9113.6]
  assign _GEN_429 = 3'h3 == _T_23937 ? shiftedStoreDataQPreg_3 : _GEN_428; // @[LoadQueue.scala 195:31:@9113.6]
  assign _GEN_430 = 3'h4 == _T_23937 ? shiftedStoreDataQPreg_4 : _GEN_429; // @[LoadQueue.scala 195:31:@9113.6]
  assign _GEN_431 = 3'h5 == _T_23937 ? shiftedStoreDataQPreg_5 : _GEN_430; // @[LoadQueue.scala 195:31:@9113.6]
  assign _GEN_432 = 3'h6 == _T_23937 ? shiftedStoreDataQPreg_6 : _GEN_431; // @[LoadQueue.scala 195:31:@9113.6]
  assign _GEN_433 = 3'h7 == _T_23937 ? shiftedStoreDataQPreg_7 : _GEN_432; // @[LoadQueue.scala 195:31:@9113.6]
  assign lastConflict_5_0 = _T_23946 ? _GEN_410 : 1'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign lastConflict_5_1 = _T_23946 ? _GEN_411 : 1'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign lastConflict_5_2 = _T_23946 ? _GEN_412 : 1'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign lastConflict_5_3 = _T_23946 ? _GEN_413 : 1'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign lastConflict_5_4 = _T_23946 ? _GEN_414 : 1'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign lastConflict_5_5 = _T_23946 ? _GEN_415 : 1'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign lastConflict_5_6 = _T_23946 ? _GEN_416 : 1'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign lastConflict_5_7 = _T_23946 ? _GEN_417 : 1'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign canBypass_5 = _T_23946 ? _GEN_425 : 1'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign bypassVal_5 = _T_23946 ? _GEN_433 : 32'h0; // @[LoadQueue.scala 192:53:@9110.4]
  assign _T_24012 = conflictPReg_6_2 ? 2'h2 : {{1'd0}, conflictPReg_6_1}; // @[LoadQueue.scala 191:60:@9143.4]
  assign _T_24013 = conflictPReg_6_3 ? 2'h3 : _T_24012; // @[LoadQueue.scala 191:60:@9144.4]
  assign _T_24014 = conflictPReg_6_4 ? 3'h4 : {{1'd0}, _T_24013}; // @[LoadQueue.scala 191:60:@9145.4]
  assign _T_24015 = conflictPReg_6_5 ? 3'h5 : _T_24014; // @[LoadQueue.scala 191:60:@9146.4]
  assign _T_24016 = conflictPReg_6_6 ? 3'h6 : _T_24015; // @[LoadQueue.scala 191:60:@9147.4]
  assign _T_24017 = conflictPReg_6_7 ? 3'h7 : _T_24016; // @[LoadQueue.scala 191:60:@9148.4]
  assign _T_24020 = conflictPReg_6_0 | conflictPReg_6_1; // @[LoadQueue.scala 192:43:@9150.4]
  assign _T_24021 = _T_24020 | conflictPReg_6_2; // @[LoadQueue.scala 192:43:@9151.4]
  assign _T_24022 = _T_24021 | conflictPReg_6_3; // @[LoadQueue.scala 192:43:@9152.4]
  assign _T_24023 = _T_24022 | conflictPReg_6_4; // @[LoadQueue.scala 192:43:@9153.4]
  assign _T_24024 = _T_24023 | conflictPReg_6_5; // @[LoadQueue.scala 192:43:@9154.4]
  assign _T_24025 = _T_24024 | conflictPReg_6_6; // @[LoadQueue.scala 192:43:@9155.4]
  assign _T_24026 = _T_24025 | conflictPReg_6_7; // @[LoadQueue.scala 192:43:@9156.4]
  assign _GEN_444 = 3'h0 == _T_24017; // @[LoadQueue.scala 193:43:@9158.6]
  assign _GEN_445 = 3'h1 == _T_24017; // @[LoadQueue.scala 193:43:@9158.6]
  assign _GEN_446 = 3'h2 == _T_24017; // @[LoadQueue.scala 193:43:@9158.6]
  assign _GEN_447 = 3'h3 == _T_24017; // @[LoadQueue.scala 193:43:@9158.6]
  assign _GEN_448 = 3'h4 == _T_24017; // @[LoadQueue.scala 193:43:@9158.6]
  assign _GEN_449 = 3'h5 == _T_24017; // @[LoadQueue.scala 193:43:@9158.6]
  assign _GEN_450 = 3'h6 == _T_24017; // @[LoadQueue.scala 193:43:@9158.6]
  assign _GEN_451 = 3'h7 == _T_24017; // @[LoadQueue.scala 193:43:@9158.6]
  assign _GEN_453 = 3'h1 == _T_24017 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@9159.6]
  assign _GEN_454 = 3'h2 == _T_24017 ? shiftedStoreDataKnownPReg_2 : _GEN_453; // @[LoadQueue.scala 194:31:@9159.6]
  assign _GEN_455 = 3'h3 == _T_24017 ? shiftedStoreDataKnownPReg_3 : _GEN_454; // @[LoadQueue.scala 194:31:@9159.6]
  assign _GEN_456 = 3'h4 == _T_24017 ? shiftedStoreDataKnownPReg_4 : _GEN_455; // @[LoadQueue.scala 194:31:@9159.6]
  assign _GEN_457 = 3'h5 == _T_24017 ? shiftedStoreDataKnownPReg_5 : _GEN_456; // @[LoadQueue.scala 194:31:@9159.6]
  assign _GEN_458 = 3'h6 == _T_24017 ? shiftedStoreDataKnownPReg_6 : _GEN_457; // @[LoadQueue.scala 194:31:@9159.6]
  assign _GEN_459 = 3'h7 == _T_24017 ? shiftedStoreDataKnownPReg_7 : _GEN_458; // @[LoadQueue.scala 194:31:@9159.6]
  assign _GEN_461 = 3'h1 == _T_24017 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@9160.6]
  assign _GEN_462 = 3'h2 == _T_24017 ? shiftedStoreDataQPreg_2 : _GEN_461; // @[LoadQueue.scala 195:31:@9160.6]
  assign _GEN_463 = 3'h3 == _T_24017 ? shiftedStoreDataQPreg_3 : _GEN_462; // @[LoadQueue.scala 195:31:@9160.6]
  assign _GEN_464 = 3'h4 == _T_24017 ? shiftedStoreDataQPreg_4 : _GEN_463; // @[LoadQueue.scala 195:31:@9160.6]
  assign _GEN_465 = 3'h5 == _T_24017 ? shiftedStoreDataQPreg_5 : _GEN_464; // @[LoadQueue.scala 195:31:@9160.6]
  assign _GEN_466 = 3'h6 == _T_24017 ? shiftedStoreDataQPreg_6 : _GEN_465; // @[LoadQueue.scala 195:31:@9160.6]
  assign _GEN_467 = 3'h7 == _T_24017 ? shiftedStoreDataQPreg_7 : _GEN_466; // @[LoadQueue.scala 195:31:@9160.6]
  assign lastConflict_6_0 = _T_24026 ? _GEN_444 : 1'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign lastConflict_6_1 = _T_24026 ? _GEN_445 : 1'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign lastConflict_6_2 = _T_24026 ? _GEN_446 : 1'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign lastConflict_6_3 = _T_24026 ? _GEN_447 : 1'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign lastConflict_6_4 = _T_24026 ? _GEN_448 : 1'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign lastConflict_6_5 = _T_24026 ? _GEN_449 : 1'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign lastConflict_6_6 = _T_24026 ? _GEN_450 : 1'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign lastConflict_6_7 = _T_24026 ? _GEN_451 : 1'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign canBypass_6 = _T_24026 ? _GEN_459 : 1'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign bypassVal_6 = _T_24026 ? _GEN_467 : 32'h0; // @[LoadQueue.scala 192:53:@9157.4]
  assign _T_24092 = conflictPReg_7_2 ? 2'h2 : {{1'd0}, conflictPReg_7_1}; // @[LoadQueue.scala 191:60:@9190.4]
  assign _T_24093 = conflictPReg_7_3 ? 2'h3 : _T_24092; // @[LoadQueue.scala 191:60:@9191.4]
  assign _T_24094 = conflictPReg_7_4 ? 3'h4 : {{1'd0}, _T_24093}; // @[LoadQueue.scala 191:60:@9192.4]
  assign _T_24095 = conflictPReg_7_5 ? 3'h5 : _T_24094; // @[LoadQueue.scala 191:60:@9193.4]
  assign _T_24096 = conflictPReg_7_6 ? 3'h6 : _T_24095; // @[LoadQueue.scala 191:60:@9194.4]
  assign _T_24097 = conflictPReg_7_7 ? 3'h7 : _T_24096; // @[LoadQueue.scala 191:60:@9195.4]
  assign _T_24100 = conflictPReg_7_0 | conflictPReg_7_1; // @[LoadQueue.scala 192:43:@9197.4]
  assign _T_24101 = _T_24100 | conflictPReg_7_2; // @[LoadQueue.scala 192:43:@9198.4]
  assign _T_24102 = _T_24101 | conflictPReg_7_3; // @[LoadQueue.scala 192:43:@9199.4]
  assign _T_24103 = _T_24102 | conflictPReg_7_4; // @[LoadQueue.scala 192:43:@9200.4]
  assign _T_24104 = _T_24103 | conflictPReg_7_5; // @[LoadQueue.scala 192:43:@9201.4]
  assign _T_24105 = _T_24104 | conflictPReg_7_6; // @[LoadQueue.scala 192:43:@9202.4]
  assign _T_24106 = _T_24105 | conflictPReg_7_7; // @[LoadQueue.scala 192:43:@9203.4]
  assign _GEN_478 = 3'h0 == _T_24097; // @[LoadQueue.scala 193:43:@9205.6]
  assign _GEN_479 = 3'h1 == _T_24097; // @[LoadQueue.scala 193:43:@9205.6]
  assign _GEN_480 = 3'h2 == _T_24097; // @[LoadQueue.scala 193:43:@9205.6]
  assign _GEN_481 = 3'h3 == _T_24097; // @[LoadQueue.scala 193:43:@9205.6]
  assign _GEN_482 = 3'h4 == _T_24097; // @[LoadQueue.scala 193:43:@9205.6]
  assign _GEN_483 = 3'h5 == _T_24097; // @[LoadQueue.scala 193:43:@9205.6]
  assign _GEN_484 = 3'h6 == _T_24097; // @[LoadQueue.scala 193:43:@9205.6]
  assign _GEN_485 = 3'h7 == _T_24097; // @[LoadQueue.scala 193:43:@9205.6]
  assign _GEN_487 = 3'h1 == _T_24097 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@9206.6]
  assign _GEN_488 = 3'h2 == _T_24097 ? shiftedStoreDataKnownPReg_2 : _GEN_487; // @[LoadQueue.scala 194:31:@9206.6]
  assign _GEN_489 = 3'h3 == _T_24097 ? shiftedStoreDataKnownPReg_3 : _GEN_488; // @[LoadQueue.scala 194:31:@9206.6]
  assign _GEN_490 = 3'h4 == _T_24097 ? shiftedStoreDataKnownPReg_4 : _GEN_489; // @[LoadQueue.scala 194:31:@9206.6]
  assign _GEN_491 = 3'h5 == _T_24097 ? shiftedStoreDataKnownPReg_5 : _GEN_490; // @[LoadQueue.scala 194:31:@9206.6]
  assign _GEN_492 = 3'h6 == _T_24097 ? shiftedStoreDataKnownPReg_6 : _GEN_491; // @[LoadQueue.scala 194:31:@9206.6]
  assign _GEN_493 = 3'h7 == _T_24097 ? shiftedStoreDataKnownPReg_7 : _GEN_492; // @[LoadQueue.scala 194:31:@9206.6]
  assign _GEN_495 = 3'h1 == _T_24097 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@9207.6]
  assign _GEN_496 = 3'h2 == _T_24097 ? shiftedStoreDataQPreg_2 : _GEN_495; // @[LoadQueue.scala 195:31:@9207.6]
  assign _GEN_497 = 3'h3 == _T_24097 ? shiftedStoreDataQPreg_3 : _GEN_496; // @[LoadQueue.scala 195:31:@9207.6]
  assign _GEN_498 = 3'h4 == _T_24097 ? shiftedStoreDataQPreg_4 : _GEN_497; // @[LoadQueue.scala 195:31:@9207.6]
  assign _GEN_499 = 3'h5 == _T_24097 ? shiftedStoreDataQPreg_5 : _GEN_498; // @[LoadQueue.scala 195:31:@9207.6]
  assign _GEN_500 = 3'h6 == _T_24097 ? shiftedStoreDataQPreg_6 : _GEN_499; // @[LoadQueue.scala 195:31:@9207.6]
  assign _GEN_501 = 3'h7 == _T_24097 ? shiftedStoreDataQPreg_7 : _GEN_500; // @[LoadQueue.scala 195:31:@9207.6]
  assign lastConflict_7_0 = _T_24106 ? _GEN_478 : 1'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign lastConflict_7_1 = _T_24106 ? _GEN_479 : 1'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign lastConflict_7_2 = _T_24106 ? _GEN_480 : 1'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign lastConflict_7_3 = _T_24106 ? _GEN_481 : 1'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign lastConflict_7_4 = _T_24106 ? _GEN_482 : 1'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign lastConflict_7_5 = _T_24106 ? _GEN_483 : 1'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign lastConflict_7_6 = _T_24106 ? _GEN_484 : 1'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign lastConflict_7_7 = _T_24106 ? _GEN_485 : 1'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign canBypass_7 = _T_24106 ? _GEN_493 : 1'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign bypassVal_7 = _T_24106 ? _GEN_501 : 32'h0; // @[LoadQueue.scala 192:53:@9204.4]
  assign _T_24150 = 8'h1 << head; // @[OneHot.scala 52:12:@9212.4]
  assign _T_24152 = _T_24150[0]; // @[util.scala 33:60:@9214.4]
  assign _T_24153 = _T_24150[1]; // @[util.scala 33:60:@9215.4]
  assign _T_24154 = _T_24150[2]; // @[util.scala 33:60:@9216.4]
  assign _T_24155 = _T_24150[3]; // @[util.scala 33:60:@9217.4]
  assign _T_24156 = _T_24150[4]; // @[util.scala 33:60:@9218.4]
  assign _T_24157 = _T_24150[5]; // @[util.scala 33:60:@9219.4]
  assign _T_24158 = _T_24150[6]; // @[util.scala 33:60:@9220.4]
  assign _T_24159 = _T_24150[7]; // @[util.scala 33:60:@9221.4]
  assign _T_25144 = dataKnownPReg_7 == 1'h0; // @[LoadQueue.scala 229:41:@9968.4]
  assign _T_25145 = addrKnownPReg_7 & _T_25144; // @[LoadQueue.scala 229:38:@9969.4]
  assign _T_25147 = bypassInitiated_7 == 1'h0; // @[LoadQueue.scala 230:12:@9971.6]
  assign _T_25149 = prevPriorityRequest_7 == 1'h0; // @[LoadQueue.scala 230:46:@9972.6]
  assign _T_25150 = _T_25147 & _T_25149; // @[LoadQueue.scala 230:43:@9973.6]
  assign _T_25152 = dataKnown_7 == 1'h0; // @[LoadQueue.scala 230:84:@9974.6]
  assign _T_25153 = _T_25150 & _T_25152; // @[LoadQueue.scala 230:81:@9975.6]
  assign _T_25156 = storeAddrNotKnownFlagsPReg_7_0 | storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 233:86:@9978.8]
  assign _T_25157 = _T_25156 | storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 233:86:@9979.8]
  assign _T_25158 = _T_25157 | storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 233:86:@9980.8]
  assign _T_25159 = _T_25158 | storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 233:86:@9981.8]
  assign _T_25160 = _T_25159 | storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 233:86:@9982.8]
  assign _T_25161 = _T_25160 | storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 233:86:@9983.8]
  assign _T_25162 = _T_25161 | storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 233:86:@9984.8]
  assign _T_25164 = _T_25162 == 1'h0; // @[LoadQueue.scala 233:38:@9985.8]
  assign _T_25175 = _T_24106 == 1'h0; // @[LoadQueue.scala 234:11:@9994.8]
  assign _T_25176 = _T_25164 & _T_25175; // @[LoadQueue.scala 233:103:@9995.8]
  assign _GEN_564 = _T_25153 ? _T_25176 : 1'h0; // @[LoadQueue.scala 230:110:@9976.6]
  assign loadRequest_7 = _T_25145 ? _GEN_564 : 1'h0; // @[LoadQueue.scala 229:71:@9970.4]
  assign _T_24184 = loadRequest_7 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9231.4]
  assign _T_25092 = dataKnownPReg_6 == 1'h0; // @[LoadQueue.scala 229:41:@9918.4]
  assign _T_25093 = addrKnownPReg_6 & _T_25092; // @[LoadQueue.scala 229:38:@9919.4]
  assign _T_25095 = bypassInitiated_6 == 1'h0; // @[LoadQueue.scala 230:12:@9921.6]
  assign _T_25097 = prevPriorityRequest_6 == 1'h0; // @[LoadQueue.scala 230:46:@9922.6]
  assign _T_25098 = _T_25095 & _T_25097; // @[LoadQueue.scala 230:43:@9923.6]
  assign _T_25100 = dataKnown_6 == 1'h0; // @[LoadQueue.scala 230:84:@9924.6]
  assign _T_25101 = _T_25098 & _T_25100; // @[LoadQueue.scala 230:81:@9925.6]
  assign _T_25104 = storeAddrNotKnownFlagsPReg_6_0 | storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 233:86:@9928.8]
  assign _T_25105 = _T_25104 | storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 233:86:@9929.8]
  assign _T_25106 = _T_25105 | storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 233:86:@9930.8]
  assign _T_25107 = _T_25106 | storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 233:86:@9931.8]
  assign _T_25108 = _T_25107 | storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 233:86:@9932.8]
  assign _T_25109 = _T_25108 | storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 233:86:@9933.8]
  assign _T_25110 = _T_25109 | storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 233:86:@9934.8]
  assign _T_25112 = _T_25110 == 1'h0; // @[LoadQueue.scala 233:38:@9935.8]
  assign _T_25123 = _T_24026 == 1'h0; // @[LoadQueue.scala 234:11:@9944.8]
  assign _T_25124 = _T_25112 & _T_25123; // @[LoadQueue.scala 233:103:@9945.8]
  assign _GEN_560 = _T_25101 ? _T_25124 : 1'h0; // @[LoadQueue.scala 230:110:@9926.6]
  assign loadRequest_6 = _T_25093 ? _GEN_560 : 1'h0; // @[LoadQueue.scala 229:71:@9920.4]
  assign _T_24185 = loadRequest_6 ? 8'h40 : _T_24184; // @[Mux.scala 31:69:@9232.4]
  assign _T_25040 = dataKnownPReg_5 == 1'h0; // @[LoadQueue.scala 229:41:@9868.4]
  assign _T_25041 = addrKnownPReg_5 & _T_25040; // @[LoadQueue.scala 229:38:@9869.4]
  assign _T_25043 = bypassInitiated_5 == 1'h0; // @[LoadQueue.scala 230:12:@9871.6]
  assign _T_25045 = prevPriorityRequest_5 == 1'h0; // @[LoadQueue.scala 230:46:@9872.6]
  assign _T_25046 = _T_25043 & _T_25045; // @[LoadQueue.scala 230:43:@9873.6]
  assign _T_25048 = dataKnown_5 == 1'h0; // @[LoadQueue.scala 230:84:@9874.6]
  assign _T_25049 = _T_25046 & _T_25048; // @[LoadQueue.scala 230:81:@9875.6]
  assign _T_25052 = storeAddrNotKnownFlagsPReg_5_0 | storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 233:86:@9878.8]
  assign _T_25053 = _T_25052 | storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 233:86:@9879.8]
  assign _T_25054 = _T_25053 | storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 233:86:@9880.8]
  assign _T_25055 = _T_25054 | storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 233:86:@9881.8]
  assign _T_25056 = _T_25055 | storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 233:86:@9882.8]
  assign _T_25057 = _T_25056 | storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 233:86:@9883.8]
  assign _T_25058 = _T_25057 | storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 233:86:@9884.8]
  assign _T_25060 = _T_25058 == 1'h0; // @[LoadQueue.scala 233:38:@9885.8]
  assign _T_25071 = _T_23946 == 1'h0; // @[LoadQueue.scala 234:11:@9894.8]
  assign _T_25072 = _T_25060 & _T_25071; // @[LoadQueue.scala 233:103:@9895.8]
  assign _GEN_556 = _T_25049 ? _T_25072 : 1'h0; // @[LoadQueue.scala 230:110:@9876.6]
  assign loadRequest_5 = _T_25041 ? _GEN_556 : 1'h0; // @[LoadQueue.scala 229:71:@9870.4]
  assign _T_24186 = loadRequest_5 ? 8'h20 : _T_24185; // @[Mux.scala 31:69:@9233.4]
  assign _T_24988 = dataKnownPReg_4 == 1'h0; // @[LoadQueue.scala 229:41:@9818.4]
  assign _T_24989 = addrKnownPReg_4 & _T_24988; // @[LoadQueue.scala 229:38:@9819.4]
  assign _T_24991 = bypassInitiated_4 == 1'h0; // @[LoadQueue.scala 230:12:@9821.6]
  assign _T_24993 = prevPriorityRequest_4 == 1'h0; // @[LoadQueue.scala 230:46:@9822.6]
  assign _T_24994 = _T_24991 & _T_24993; // @[LoadQueue.scala 230:43:@9823.6]
  assign _T_24996 = dataKnown_4 == 1'h0; // @[LoadQueue.scala 230:84:@9824.6]
  assign _T_24997 = _T_24994 & _T_24996; // @[LoadQueue.scala 230:81:@9825.6]
  assign _T_25000 = storeAddrNotKnownFlagsPReg_4_0 | storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 233:86:@9828.8]
  assign _T_25001 = _T_25000 | storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 233:86:@9829.8]
  assign _T_25002 = _T_25001 | storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 233:86:@9830.8]
  assign _T_25003 = _T_25002 | storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 233:86:@9831.8]
  assign _T_25004 = _T_25003 | storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 233:86:@9832.8]
  assign _T_25005 = _T_25004 | storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 233:86:@9833.8]
  assign _T_25006 = _T_25005 | storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 233:86:@9834.8]
  assign _T_25008 = _T_25006 == 1'h0; // @[LoadQueue.scala 233:38:@9835.8]
  assign _T_25019 = _T_23866 == 1'h0; // @[LoadQueue.scala 234:11:@9844.8]
  assign _T_25020 = _T_25008 & _T_25019; // @[LoadQueue.scala 233:103:@9845.8]
  assign _GEN_552 = _T_24997 ? _T_25020 : 1'h0; // @[LoadQueue.scala 230:110:@9826.6]
  assign loadRequest_4 = _T_24989 ? _GEN_552 : 1'h0; // @[LoadQueue.scala 229:71:@9820.4]
  assign _T_24187 = loadRequest_4 ? 8'h10 : _T_24186; // @[Mux.scala 31:69:@9234.4]
  assign _T_24936 = dataKnownPReg_3 == 1'h0; // @[LoadQueue.scala 229:41:@9768.4]
  assign _T_24937 = addrKnownPReg_3 & _T_24936; // @[LoadQueue.scala 229:38:@9769.4]
  assign _T_24939 = bypassInitiated_3 == 1'h0; // @[LoadQueue.scala 230:12:@9771.6]
  assign _T_24941 = prevPriorityRequest_3 == 1'h0; // @[LoadQueue.scala 230:46:@9772.6]
  assign _T_24942 = _T_24939 & _T_24941; // @[LoadQueue.scala 230:43:@9773.6]
  assign _T_24944 = dataKnown_3 == 1'h0; // @[LoadQueue.scala 230:84:@9774.6]
  assign _T_24945 = _T_24942 & _T_24944; // @[LoadQueue.scala 230:81:@9775.6]
  assign _T_24948 = storeAddrNotKnownFlagsPReg_3_0 | storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 233:86:@9778.8]
  assign _T_24949 = _T_24948 | storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 233:86:@9779.8]
  assign _T_24950 = _T_24949 | storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 233:86:@9780.8]
  assign _T_24951 = _T_24950 | storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 233:86:@9781.8]
  assign _T_24952 = _T_24951 | storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 233:86:@9782.8]
  assign _T_24953 = _T_24952 | storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 233:86:@9783.8]
  assign _T_24954 = _T_24953 | storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 233:86:@9784.8]
  assign _T_24956 = _T_24954 == 1'h0; // @[LoadQueue.scala 233:38:@9785.8]
  assign _T_24967 = _T_23786 == 1'h0; // @[LoadQueue.scala 234:11:@9794.8]
  assign _T_24968 = _T_24956 & _T_24967; // @[LoadQueue.scala 233:103:@9795.8]
  assign _GEN_548 = _T_24945 ? _T_24968 : 1'h0; // @[LoadQueue.scala 230:110:@9776.6]
  assign loadRequest_3 = _T_24937 ? _GEN_548 : 1'h0; // @[LoadQueue.scala 229:71:@9770.4]
  assign _T_24188 = loadRequest_3 ? 8'h8 : _T_24187; // @[Mux.scala 31:69:@9235.4]
  assign _T_24884 = dataKnownPReg_2 == 1'h0; // @[LoadQueue.scala 229:41:@9718.4]
  assign _T_24885 = addrKnownPReg_2 & _T_24884; // @[LoadQueue.scala 229:38:@9719.4]
  assign _T_24887 = bypassInitiated_2 == 1'h0; // @[LoadQueue.scala 230:12:@9721.6]
  assign _T_24889 = prevPriorityRequest_2 == 1'h0; // @[LoadQueue.scala 230:46:@9722.6]
  assign _T_24890 = _T_24887 & _T_24889; // @[LoadQueue.scala 230:43:@9723.6]
  assign _T_24892 = dataKnown_2 == 1'h0; // @[LoadQueue.scala 230:84:@9724.6]
  assign _T_24893 = _T_24890 & _T_24892; // @[LoadQueue.scala 230:81:@9725.6]
  assign _T_24896 = storeAddrNotKnownFlagsPReg_2_0 | storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 233:86:@9728.8]
  assign _T_24897 = _T_24896 | storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 233:86:@9729.8]
  assign _T_24898 = _T_24897 | storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 233:86:@9730.8]
  assign _T_24899 = _T_24898 | storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 233:86:@9731.8]
  assign _T_24900 = _T_24899 | storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 233:86:@9732.8]
  assign _T_24901 = _T_24900 | storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 233:86:@9733.8]
  assign _T_24902 = _T_24901 | storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 233:86:@9734.8]
  assign _T_24904 = _T_24902 == 1'h0; // @[LoadQueue.scala 233:38:@9735.8]
  assign _T_24915 = _T_23706 == 1'h0; // @[LoadQueue.scala 234:11:@9744.8]
  assign _T_24916 = _T_24904 & _T_24915; // @[LoadQueue.scala 233:103:@9745.8]
  assign _GEN_544 = _T_24893 ? _T_24916 : 1'h0; // @[LoadQueue.scala 230:110:@9726.6]
  assign loadRequest_2 = _T_24885 ? _GEN_544 : 1'h0; // @[LoadQueue.scala 229:71:@9720.4]
  assign _T_24189 = loadRequest_2 ? 8'h4 : _T_24188; // @[Mux.scala 31:69:@9236.4]
  assign _T_24832 = dataKnownPReg_1 == 1'h0; // @[LoadQueue.scala 229:41:@9668.4]
  assign _T_24833 = addrKnownPReg_1 & _T_24832; // @[LoadQueue.scala 229:38:@9669.4]
  assign _T_24835 = bypassInitiated_1 == 1'h0; // @[LoadQueue.scala 230:12:@9671.6]
  assign _T_24837 = prevPriorityRequest_1 == 1'h0; // @[LoadQueue.scala 230:46:@9672.6]
  assign _T_24838 = _T_24835 & _T_24837; // @[LoadQueue.scala 230:43:@9673.6]
  assign _T_24840 = dataKnown_1 == 1'h0; // @[LoadQueue.scala 230:84:@9674.6]
  assign _T_24841 = _T_24838 & _T_24840; // @[LoadQueue.scala 230:81:@9675.6]
  assign _T_24844 = storeAddrNotKnownFlagsPReg_1_0 | storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 233:86:@9678.8]
  assign _T_24845 = _T_24844 | storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 233:86:@9679.8]
  assign _T_24846 = _T_24845 | storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 233:86:@9680.8]
  assign _T_24847 = _T_24846 | storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 233:86:@9681.8]
  assign _T_24848 = _T_24847 | storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 233:86:@9682.8]
  assign _T_24849 = _T_24848 | storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 233:86:@9683.8]
  assign _T_24850 = _T_24849 | storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 233:86:@9684.8]
  assign _T_24852 = _T_24850 == 1'h0; // @[LoadQueue.scala 233:38:@9685.8]
  assign _T_24863 = _T_23626 == 1'h0; // @[LoadQueue.scala 234:11:@9694.8]
  assign _T_24864 = _T_24852 & _T_24863; // @[LoadQueue.scala 233:103:@9695.8]
  assign _GEN_540 = _T_24841 ? _T_24864 : 1'h0; // @[LoadQueue.scala 230:110:@9676.6]
  assign loadRequest_1 = _T_24833 ? _GEN_540 : 1'h0; // @[LoadQueue.scala 229:71:@9670.4]
  assign _T_24190 = loadRequest_1 ? 8'h2 : _T_24189; // @[Mux.scala 31:69:@9237.4]
  assign _T_24780 = dataKnownPReg_0 == 1'h0; // @[LoadQueue.scala 229:41:@9618.4]
  assign _T_24781 = addrKnownPReg_0 & _T_24780; // @[LoadQueue.scala 229:38:@9619.4]
  assign _T_24783 = bypassInitiated_0 == 1'h0; // @[LoadQueue.scala 230:12:@9621.6]
  assign _T_24785 = prevPriorityRequest_0 == 1'h0; // @[LoadQueue.scala 230:46:@9622.6]
  assign _T_24786 = _T_24783 & _T_24785; // @[LoadQueue.scala 230:43:@9623.6]
  assign _T_24788 = dataKnown_0 == 1'h0; // @[LoadQueue.scala 230:84:@9624.6]
  assign _T_24789 = _T_24786 & _T_24788; // @[LoadQueue.scala 230:81:@9625.6]
  assign _T_24792 = storeAddrNotKnownFlagsPReg_0_0 | storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 233:86:@9628.8]
  assign _T_24793 = _T_24792 | storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 233:86:@9629.8]
  assign _T_24794 = _T_24793 | storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 233:86:@9630.8]
  assign _T_24795 = _T_24794 | storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 233:86:@9631.8]
  assign _T_24796 = _T_24795 | storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 233:86:@9632.8]
  assign _T_24797 = _T_24796 | storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 233:86:@9633.8]
  assign _T_24798 = _T_24797 | storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 233:86:@9634.8]
  assign _T_24800 = _T_24798 == 1'h0; // @[LoadQueue.scala 233:38:@9635.8]
  assign _T_24811 = _T_23546 == 1'h0; // @[LoadQueue.scala 234:11:@9644.8]
  assign _T_24812 = _T_24800 & _T_24811; // @[LoadQueue.scala 233:103:@9645.8]
  assign _GEN_536 = _T_24789 ? _T_24812 : 1'h0; // @[LoadQueue.scala 230:110:@9626.6]
  assign loadRequest_0 = _T_24781 ? _GEN_536 : 1'h0; // @[LoadQueue.scala 229:71:@9620.4]
  assign _T_24191 = loadRequest_0 ? 8'h1 : _T_24190; // @[Mux.scala 31:69:@9238.4]
  assign _T_24192 = _T_24191[0]; // @[OneHot.scala 66:30:@9239.4]
  assign _T_24193 = _T_24191[1]; // @[OneHot.scala 66:30:@9240.4]
  assign _T_24194 = _T_24191[2]; // @[OneHot.scala 66:30:@9241.4]
  assign _T_24195 = _T_24191[3]; // @[OneHot.scala 66:30:@9242.4]
  assign _T_24196 = _T_24191[4]; // @[OneHot.scala 66:30:@9243.4]
  assign _T_24197 = _T_24191[5]; // @[OneHot.scala 66:30:@9244.4]
  assign _T_24198 = _T_24191[6]; // @[OneHot.scala 66:30:@9245.4]
  assign _T_24199 = _T_24191[7]; // @[OneHot.scala 66:30:@9246.4]
  assign _T_24224 = loadRequest_0 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9256.4]
  assign _T_24225 = loadRequest_7 ? 8'h40 : _T_24224; // @[Mux.scala 31:69:@9257.4]
  assign _T_24226 = loadRequest_6 ? 8'h20 : _T_24225; // @[Mux.scala 31:69:@9258.4]
  assign _T_24227 = loadRequest_5 ? 8'h10 : _T_24226; // @[Mux.scala 31:69:@9259.4]
  assign _T_24228 = loadRequest_4 ? 8'h8 : _T_24227; // @[Mux.scala 31:69:@9260.4]
  assign _T_24229 = loadRequest_3 ? 8'h4 : _T_24228; // @[Mux.scala 31:69:@9261.4]
  assign _T_24230 = loadRequest_2 ? 8'h2 : _T_24229; // @[Mux.scala 31:69:@9262.4]
  assign _T_24231 = loadRequest_1 ? 8'h1 : _T_24230; // @[Mux.scala 31:69:@9263.4]
  assign _T_24232 = _T_24231[0]; // @[OneHot.scala 66:30:@9264.4]
  assign _T_24233 = _T_24231[1]; // @[OneHot.scala 66:30:@9265.4]
  assign _T_24234 = _T_24231[2]; // @[OneHot.scala 66:30:@9266.4]
  assign _T_24235 = _T_24231[3]; // @[OneHot.scala 66:30:@9267.4]
  assign _T_24236 = _T_24231[4]; // @[OneHot.scala 66:30:@9268.4]
  assign _T_24237 = _T_24231[5]; // @[OneHot.scala 66:30:@9269.4]
  assign _T_24238 = _T_24231[6]; // @[OneHot.scala 66:30:@9270.4]
  assign _T_24239 = _T_24231[7]; // @[OneHot.scala 66:30:@9271.4]
  assign _T_24264 = loadRequest_1 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9281.4]
  assign _T_24265 = loadRequest_0 ? 8'h40 : _T_24264; // @[Mux.scala 31:69:@9282.4]
  assign _T_24266 = loadRequest_7 ? 8'h20 : _T_24265; // @[Mux.scala 31:69:@9283.4]
  assign _T_24267 = loadRequest_6 ? 8'h10 : _T_24266; // @[Mux.scala 31:69:@9284.4]
  assign _T_24268 = loadRequest_5 ? 8'h8 : _T_24267; // @[Mux.scala 31:69:@9285.4]
  assign _T_24269 = loadRequest_4 ? 8'h4 : _T_24268; // @[Mux.scala 31:69:@9286.4]
  assign _T_24270 = loadRequest_3 ? 8'h2 : _T_24269; // @[Mux.scala 31:69:@9287.4]
  assign _T_24271 = loadRequest_2 ? 8'h1 : _T_24270; // @[Mux.scala 31:69:@9288.4]
  assign _T_24272 = _T_24271[0]; // @[OneHot.scala 66:30:@9289.4]
  assign _T_24273 = _T_24271[1]; // @[OneHot.scala 66:30:@9290.4]
  assign _T_24274 = _T_24271[2]; // @[OneHot.scala 66:30:@9291.4]
  assign _T_24275 = _T_24271[3]; // @[OneHot.scala 66:30:@9292.4]
  assign _T_24276 = _T_24271[4]; // @[OneHot.scala 66:30:@9293.4]
  assign _T_24277 = _T_24271[5]; // @[OneHot.scala 66:30:@9294.4]
  assign _T_24278 = _T_24271[6]; // @[OneHot.scala 66:30:@9295.4]
  assign _T_24279 = _T_24271[7]; // @[OneHot.scala 66:30:@9296.4]
  assign _T_24304 = loadRequest_2 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9306.4]
  assign _T_24305 = loadRequest_1 ? 8'h40 : _T_24304; // @[Mux.scala 31:69:@9307.4]
  assign _T_24306 = loadRequest_0 ? 8'h20 : _T_24305; // @[Mux.scala 31:69:@9308.4]
  assign _T_24307 = loadRequest_7 ? 8'h10 : _T_24306; // @[Mux.scala 31:69:@9309.4]
  assign _T_24308 = loadRequest_6 ? 8'h8 : _T_24307; // @[Mux.scala 31:69:@9310.4]
  assign _T_24309 = loadRequest_5 ? 8'h4 : _T_24308; // @[Mux.scala 31:69:@9311.4]
  assign _T_24310 = loadRequest_4 ? 8'h2 : _T_24309; // @[Mux.scala 31:69:@9312.4]
  assign _T_24311 = loadRequest_3 ? 8'h1 : _T_24310; // @[Mux.scala 31:69:@9313.4]
  assign _T_24312 = _T_24311[0]; // @[OneHot.scala 66:30:@9314.4]
  assign _T_24313 = _T_24311[1]; // @[OneHot.scala 66:30:@9315.4]
  assign _T_24314 = _T_24311[2]; // @[OneHot.scala 66:30:@9316.4]
  assign _T_24315 = _T_24311[3]; // @[OneHot.scala 66:30:@9317.4]
  assign _T_24316 = _T_24311[4]; // @[OneHot.scala 66:30:@9318.4]
  assign _T_24317 = _T_24311[5]; // @[OneHot.scala 66:30:@9319.4]
  assign _T_24318 = _T_24311[6]; // @[OneHot.scala 66:30:@9320.4]
  assign _T_24319 = _T_24311[7]; // @[OneHot.scala 66:30:@9321.4]
  assign _T_24344 = loadRequest_3 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9331.4]
  assign _T_24345 = loadRequest_2 ? 8'h40 : _T_24344; // @[Mux.scala 31:69:@9332.4]
  assign _T_24346 = loadRequest_1 ? 8'h20 : _T_24345; // @[Mux.scala 31:69:@9333.4]
  assign _T_24347 = loadRequest_0 ? 8'h10 : _T_24346; // @[Mux.scala 31:69:@9334.4]
  assign _T_24348 = loadRequest_7 ? 8'h8 : _T_24347; // @[Mux.scala 31:69:@9335.4]
  assign _T_24349 = loadRequest_6 ? 8'h4 : _T_24348; // @[Mux.scala 31:69:@9336.4]
  assign _T_24350 = loadRequest_5 ? 8'h2 : _T_24349; // @[Mux.scala 31:69:@9337.4]
  assign _T_24351 = loadRequest_4 ? 8'h1 : _T_24350; // @[Mux.scala 31:69:@9338.4]
  assign _T_24352 = _T_24351[0]; // @[OneHot.scala 66:30:@9339.4]
  assign _T_24353 = _T_24351[1]; // @[OneHot.scala 66:30:@9340.4]
  assign _T_24354 = _T_24351[2]; // @[OneHot.scala 66:30:@9341.4]
  assign _T_24355 = _T_24351[3]; // @[OneHot.scala 66:30:@9342.4]
  assign _T_24356 = _T_24351[4]; // @[OneHot.scala 66:30:@9343.4]
  assign _T_24357 = _T_24351[5]; // @[OneHot.scala 66:30:@9344.4]
  assign _T_24358 = _T_24351[6]; // @[OneHot.scala 66:30:@9345.4]
  assign _T_24359 = _T_24351[7]; // @[OneHot.scala 66:30:@9346.4]
  assign _T_24384 = loadRequest_4 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9356.4]
  assign _T_24385 = loadRequest_3 ? 8'h40 : _T_24384; // @[Mux.scala 31:69:@9357.4]
  assign _T_24386 = loadRequest_2 ? 8'h20 : _T_24385; // @[Mux.scala 31:69:@9358.4]
  assign _T_24387 = loadRequest_1 ? 8'h10 : _T_24386; // @[Mux.scala 31:69:@9359.4]
  assign _T_24388 = loadRequest_0 ? 8'h8 : _T_24387; // @[Mux.scala 31:69:@9360.4]
  assign _T_24389 = loadRequest_7 ? 8'h4 : _T_24388; // @[Mux.scala 31:69:@9361.4]
  assign _T_24390 = loadRequest_6 ? 8'h2 : _T_24389; // @[Mux.scala 31:69:@9362.4]
  assign _T_24391 = loadRequest_5 ? 8'h1 : _T_24390; // @[Mux.scala 31:69:@9363.4]
  assign _T_24392 = _T_24391[0]; // @[OneHot.scala 66:30:@9364.4]
  assign _T_24393 = _T_24391[1]; // @[OneHot.scala 66:30:@9365.4]
  assign _T_24394 = _T_24391[2]; // @[OneHot.scala 66:30:@9366.4]
  assign _T_24395 = _T_24391[3]; // @[OneHot.scala 66:30:@9367.4]
  assign _T_24396 = _T_24391[4]; // @[OneHot.scala 66:30:@9368.4]
  assign _T_24397 = _T_24391[5]; // @[OneHot.scala 66:30:@9369.4]
  assign _T_24398 = _T_24391[6]; // @[OneHot.scala 66:30:@9370.4]
  assign _T_24399 = _T_24391[7]; // @[OneHot.scala 66:30:@9371.4]
  assign _T_24424 = loadRequest_5 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9381.4]
  assign _T_24425 = loadRequest_4 ? 8'h40 : _T_24424; // @[Mux.scala 31:69:@9382.4]
  assign _T_24426 = loadRequest_3 ? 8'h20 : _T_24425; // @[Mux.scala 31:69:@9383.4]
  assign _T_24427 = loadRequest_2 ? 8'h10 : _T_24426; // @[Mux.scala 31:69:@9384.4]
  assign _T_24428 = loadRequest_1 ? 8'h8 : _T_24427; // @[Mux.scala 31:69:@9385.4]
  assign _T_24429 = loadRequest_0 ? 8'h4 : _T_24428; // @[Mux.scala 31:69:@9386.4]
  assign _T_24430 = loadRequest_7 ? 8'h2 : _T_24429; // @[Mux.scala 31:69:@9387.4]
  assign _T_24431 = loadRequest_6 ? 8'h1 : _T_24430; // @[Mux.scala 31:69:@9388.4]
  assign _T_24432 = _T_24431[0]; // @[OneHot.scala 66:30:@9389.4]
  assign _T_24433 = _T_24431[1]; // @[OneHot.scala 66:30:@9390.4]
  assign _T_24434 = _T_24431[2]; // @[OneHot.scala 66:30:@9391.4]
  assign _T_24435 = _T_24431[3]; // @[OneHot.scala 66:30:@9392.4]
  assign _T_24436 = _T_24431[4]; // @[OneHot.scala 66:30:@9393.4]
  assign _T_24437 = _T_24431[5]; // @[OneHot.scala 66:30:@9394.4]
  assign _T_24438 = _T_24431[6]; // @[OneHot.scala 66:30:@9395.4]
  assign _T_24439 = _T_24431[7]; // @[OneHot.scala 66:30:@9396.4]
  assign _T_24464 = loadRequest_6 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@9406.4]
  assign _T_24465 = loadRequest_5 ? 8'h40 : _T_24464; // @[Mux.scala 31:69:@9407.4]
  assign _T_24466 = loadRequest_4 ? 8'h20 : _T_24465; // @[Mux.scala 31:69:@9408.4]
  assign _T_24467 = loadRequest_3 ? 8'h10 : _T_24466; // @[Mux.scala 31:69:@9409.4]
  assign _T_24468 = loadRequest_2 ? 8'h8 : _T_24467; // @[Mux.scala 31:69:@9410.4]
  assign _T_24469 = loadRequest_1 ? 8'h4 : _T_24468; // @[Mux.scala 31:69:@9411.4]
  assign _T_24470 = loadRequest_0 ? 8'h2 : _T_24469; // @[Mux.scala 31:69:@9412.4]
  assign _T_24471 = loadRequest_7 ? 8'h1 : _T_24470; // @[Mux.scala 31:69:@9413.4]
  assign _T_24472 = _T_24471[0]; // @[OneHot.scala 66:30:@9414.4]
  assign _T_24473 = _T_24471[1]; // @[OneHot.scala 66:30:@9415.4]
  assign _T_24474 = _T_24471[2]; // @[OneHot.scala 66:30:@9416.4]
  assign _T_24475 = _T_24471[3]; // @[OneHot.scala 66:30:@9417.4]
  assign _T_24476 = _T_24471[4]; // @[OneHot.scala 66:30:@9418.4]
  assign _T_24477 = _T_24471[5]; // @[OneHot.scala 66:30:@9419.4]
  assign _T_24478 = _T_24471[6]; // @[OneHot.scala 66:30:@9420.4]
  assign _T_24479 = _T_24471[7]; // @[OneHot.scala 66:30:@9421.4]
  assign _T_24520 = {_T_24199,_T_24198,_T_24197,_T_24196,_T_24195,_T_24194,_T_24193,_T_24192}; // @[Mux.scala 19:72:@9437.4]
  assign _T_24522 = _T_24152 ? _T_24520 : 8'h0; // @[Mux.scala 19:72:@9438.4]
  assign _T_24529 = {_T_24238,_T_24237,_T_24236,_T_24235,_T_24234,_T_24233,_T_24232,_T_24239}; // @[Mux.scala 19:72:@9445.4]
  assign _T_24531 = _T_24153 ? _T_24529 : 8'h0; // @[Mux.scala 19:72:@9446.4]
  assign _T_24538 = {_T_24277,_T_24276,_T_24275,_T_24274,_T_24273,_T_24272,_T_24279,_T_24278}; // @[Mux.scala 19:72:@9453.4]
  assign _T_24540 = _T_24154 ? _T_24538 : 8'h0; // @[Mux.scala 19:72:@9454.4]
  assign _T_24547 = {_T_24316,_T_24315,_T_24314,_T_24313,_T_24312,_T_24319,_T_24318,_T_24317}; // @[Mux.scala 19:72:@9461.4]
  assign _T_24549 = _T_24155 ? _T_24547 : 8'h0; // @[Mux.scala 19:72:@9462.4]
  assign _T_24556 = {_T_24355,_T_24354,_T_24353,_T_24352,_T_24359,_T_24358,_T_24357,_T_24356}; // @[Mux.scala 19:72:@9469.4]
  assign _T_24558 = _T_24156 ? _T_24556 : 8'h0; // @[Mux.scala 19:72:@9470.4]
  assign _T_24565 = {_T_24394,_T_24393,_T_24392,_T_24399,_T_24398,_T_24397,_T_24396,_T_24395}; // @[Mux.scala 19:72:@9477.4]
  assign _T_24567 = _T_24157 ? _T_24565 : 8'h0; // @[Mux.scala 19:72:@9478.4]
  assign _T_24574 = {_T_24433,_T_24432,_T_24439,_T_24438,_T_24437,_T_24436,_T_24435,_T_24434}; // @[Mux.scala 19:72:@9485.4]
  assign _T_24576 = _T_24158 ? _T_24574 : 8'h0; // @[Mux.scala 19:72:@9486.4]
  assign _T_24583 = {_T_24472,_T_24479,_T_24478,_T_24477,_T_24476,_T_24475,_T_24474,_T_24473}; // @[Mux.scala 19:72:@9493.4]
  assign _T_24585 = _T_24159 ? _T_24583 : 8'h0; // @[Mux.scala 19:72:@9494.4]
  assign _T_24586 = _T_24522 | _T_24531; // @[Mux.scala 19:72:@9495.4]
  assign _T_24587 = _T_24586 | _T_24540; // @[Mux.scala 19:72:@9496.4]
  assign _T_24588 = _T_24587 | _T_24549; // @[Mux.scala 19:72:@9497.4]
  assign _T_24589 = _T_24588 | _T_24558; // @[Mux.scala 19:72:@9498.4]
  assign _T_24590 = _T_24589 | _T_24567; // @[Mux.scala 19:72:@9499.4]
  assign _T_24591 = _T_24590 | _T_24576; // @[Mux.scala 19:72:@9500.4]
  assign _T_24592 = _T_24591 | _T_24585; // @[Mux.scala 19:72:@9501.4]
  assign priorityLoadRequest_0 = _T_24592[0]; // @[Mux.scala 19:72:@9505.4]
  assign priorityLoadRequest_1 = _T_24592[1]; // @[Mux.scala 19:72:@9507.4]
  assign priorityLoadRequest_2 = _T_24592[2]; // @[Mux.scala 19:72:@9509.4]
  assign priorityLoadRequest_3 = _T_24592[3]; // @[Mux.scala 19:72:@9511.4]
  assign priorityLoadRequest_4 = _T_24592[4]; // @[Mux.scala 19:72:@9513.4]
  assign priorityLoadRequest_5 = _T_24592[5]; // @[Mux.scala 19:72:@9515.4]
  assign priorityLoadRequest_6 = _T_24592[6]; // @[Mux.scala 19:72:@9517.4]
  assign priorityLoadRequest_7 = _T_24592[7]; // @[Mux.scala 19:72:@9519.4]
  assign _GEN_512 = io_memIsReadyForLoads ? priorityLoadRequest_0 : 1'h0; // @[LoadQueue.scala 208:31:@9531.4]
  assign _GEN_513 = io_memIsReadyForLoads ? priorityLoadRequest_1 : 1'h0; // @[LoadQueue.scala 208:31:@9531.4]
  assign _GEN_514 = io_memIsReadyForLoads ? priorityLoadRequest_2 : 1'h0; // @[LoadQueue.scala 208:31:@9531.4]
  assign _GEN_515 = io_memIsReadyForLoads ? priorityLoadRequest_3 : 1'h0; // @[LoadQueue.scala 208:31:@9531.4]
  assign _GEN_516 = io_memIsReadyForLoads ? priorityLoadRequest_4 : 1'h0; // @[LoadQueue.scala 208:31:@9531.4]
  assign _GEN_517 = io_memIsReadyForLoads ? priorityLoadRequest_5 : 1'h0; // @[LoadQueue.scala 208:31:@9531.4]
  assign _GEN_518 = io_memIsReadyForLoads ? priorityLoadRequest_6 : 1'h0; // @[LoadQueue.scala 208:31:@9531.4]
  assign _GEN_519 = io_memIsReadyForLoads ? priorityLoadRequest_7 : 1'h0; // @[LoadQueue.scala 208:31:@9531.4]
  assign _T_24819 = {storeAddrNotKnownFlagsPReg_0_7,storeAddrNotKnownFlagsPReg_0_6,storeAddrNotKnownFlagsPReg_0_5,storeAddrNotKnownFlagsPReg_0_4,storeAddrNotKnownFlagsPReg_0_3,storeAddrNotKnownFlagsPReg_0_2,storeAddrNotKnownFlagsPReg_0_1,storeAddrNotKnownFlagsPReg_0_0}; // @[LoadQueue.scala 238:58:@9653.8]
  assign _T_24826 = {lastConflict_0_7,lastConflict_0_6,lastConflict_0_5,lastConflict_0_4,lastConflict_0_3,lastConflict_0_2,lastConflict_0_1,lastConflict_0_0}; // @[LoadQueue.scala 238:96:@9660.8]
  assign _T_24827 = _T_24819 < _T_24826; // @[LoadQueue.scala 238:61:@9661.8]
  assign _T_24828 = canBypass_0 & _T_24827; // @[LoadQueue.scala 237:64:@9662.8]
  assign _GEN_537 = _T_24789 ? _T_24828 : 1'h0; // @[LoadQueue.scala 230:110:@9626.6]
  assign bypassRequest_0 = _T_24781 ? _GEN_537 : 1'h0; // @[LoadQueue.scala 229:71:@9620.4]
  assign _GEN_520 = bypassRequest_0 ? 1'h1 : bypassInitiated_0; // @[LoadQueue.scala 217:34:@9564.6]
  assign _GEN_521 = initBits_0 ? 1'h0 : _GEN_520; // @[LoadQueue.scala 215:23:@9560.4]
  assign _T_24871 = {storeAddrNotKnownFlagsPReg_1_7,storeAddrNotKnownFlagsPReg_1_6,storeAddrNotKnownFlagsPReg_1_5,storeAddrNotKnownFlagsPReg_1_4,storeAddrNotKnownFlagsPReg_1_3,storeAddrNotKnownFlagsPReg_1_2,storeAddrNotKnownFlagsPReg_1_1,storeAddrNotKnownFlagsPReg_1_0}; // @[LoadQueue.scala 238:58:@9703.8]
  assign _T_24878 = {lastConflict_1_7,lastConflict_1_6,lastConflict_1_5,lastConflict_1_4,lastConflict_1_3,lastConflict_1_2,lastConflict_1_1,lastConflict_1_0}; // @[LoadQueue.scala 238:96:@9710.8]
  assign _T_24879 = _T_24871 < _T_24878; // @[LoadQueue.scala 238:61:@9711.8]
  assign _T_24880 = canBypass_1 & _T_24879; // @[LoadQueue.scala 237:64:@9712.8]
  assign _GEN_541 = _T_24841 ? _T_24880 : 1'h0; // @[LoadQueue.scala 230:110:@9676.6]
  assign bypassRequest_1 = _T_24833 ? _GEN_541 : 1'h0; // @[LoadQueue.scala 229:71:@9670.4]
  assign _GEN_522 = bypassRequest_1 ? 1'h1 : bypassInitiated_1; // @[LoadQueue.scala 217:34:@9571.6]
  assign _GEN_523 = initBits_1 ? 1'h0 : _GEN_522; // @[LoadQueue.scala 215:23:@9567.4]
  assign _T_24923 = {storeAddrNotKnownFlagsPReg_2_7,storeAddrNotKnownFlagsPReg_2_6,storeAddrNotKnownFlagsPReg_2_5,storeAddrNotKnownFlagsPReg_2_4,storeAddrNotKnownFlagsPReg_2_3,storeAddrNotKnownFlagsPReg_2_2,storeAddrNotKnownFlagsPReg_2_1,storeAddrNotKnownFlagsPReg_2_0}; // @[LoadQueue.scala 238:58:@9753.8]
  assign _T_24930 = {lastConflict_2_7,lastConflict_2_6,lastConflict_2_5,lastConflict_2_4,lastConflict_2_3,lastConflict_2_2,lastConflict_2_1,lastConflict_2_0}; // @[LoadQueue.scala 238:96:@9760.8]
  assign _T_24931 = _T_24923 < _T_24930; // @[LoadQueue.scala 238:61:@9761.8]
  assign _T_24932 = canBypass_2 & _T_24931; // @[LoadQueue.scala 237:64:@9762.8]
  assign _GEN_545 = _T_24893 ? _T_24932 : 1'h0; // @[LoadQueue.scala 230:110:@9726.6]
  assign bypassRequest_2 = _T_24885 ? _GEN_545 : 1'h0; // @[LoadQueue.scala 229:71:@9720.4]
  assign _GEN_524 = bypassRequest_2 ? 1'h1 : bypassInitiated_2; // @[LoadQueue.scala 217:34:@9578.6]
  assign _GEN_525 = initBits_2 ? 1'h0 : _GEN_524; // @[LoadQueue.scala 215:23:@9574.4]
  assign _T_24975 = {storeAddrNotKnownFlagsPReg_3_7,storeAddrNotKnownFlagsPReg_3_6,storeAddrNotKnownFlagsPReg_3_5,storeAddrNotKnownFlagsPReg_3_4,storeAddrNotKnownFlagsPReg_3_3,storeAddrNotKnownFlagsPReg_3_2,storeAddrNotKnownFlagsPReg_3_1,storeAddrNotKnownFlagsPReg_3_0}; // @[LoadQueue.scala 238:58:@9803.8]
  assign _T_24982 = {lastConflict_3_7,lastConflict_3_6,lastConflict_3_5,lastConflict_3_4,lastConflict_3_3,lastConflict_3_2,lastConflict_3_1,lastConflict_3_0}; // @[LoadQueue.scala 238:96:@9810.8]
  assign _T_24983 = _T_24975 < _T_24982; // @[LoadQueue.scala 238:61:@9811.8]
  assign _T_24984 = canBypass_3 & _T_24983; // @[LoadQueue.scala 237:64:@9812.8]
  assign _GEN_549 = _T_24945 ? _T_24984 : 1'h0; // @[LoadQueue.scala 230:110:@9776.6]
  assign bypassRequest_3 = _T_24937 ? _GEN_549 : 1'h0; // @[LoadQueue.scala 229:71:@9770.4]
  assign _GEN_526 = bypassRequest_3 ? 1'h1 : bypassInitiated_3; // @[LoadQueue.scala 217:34:@9585.6]
  assign _GEN_527 = initBits_3 ? 1'h0 : _GEN_526; // @[LoadQueue.scala 215:23:@9581.4]
  assign _T_25027 = {storeAddrNotKnownFlagsPReg_4_7,storeAddrNotKnownFlagsPReg_4_6,storeAddrNotKnownFlagsPReg_4_5,storeAddrNotKnownFlagsPReg_4_4,storeAddrNotKnownFlagsPReg_4_3,storeAddrNotKnownFlagsPReg_4_2,storeAddrNotKnownFlagsPReg_4_1,storeAddrNotKnownFlagsPReg_4_0}; // @[LoadQueue.scala 238:58:@9853.8]
  assign _T_25034 = {lastConflict_4_7,lastConflict_4_6,lastConflict_4_5,lastConflict_4_4,lastConflict_4_3,lastConflict_4_2,lastConflict_4_1,lastConflict_4_0}; // @[LoadQueue.scala 238:96:@9860.8]
  assign _T_25035 = _T_25027 < _T_25034; // @[LoadQueue.scala 238:61:@9861.8]
  assign _T_25036 = canBypass_4 & _T_25035; // @[LoadQueue.scala 237:64:@9862.8]
  assign _GEN_553 = _T_24997 ? _T_25036 : 1'h0; // @[LoadQueue.scala 230:110:@9826.6]
  assign bypassRequest_4 = _T_24989 ? _GEN_553 : 1'h0; // @[LoadQueue.scala 229:71:@9820.4]
  assign _GEN_528 = bypassRequest_4 ? 1'h1 : bypassInitiated_4; // @[LoadQueue.scala 217:34:@9592.6]
  assign _GEN_529 = initBits_4 ? 1'h0 : _GEN_528; // @[LoadQueue.scala 215:23:@9588.4]
  assign _T_25079 = {storeAddrNotKnownFlagsPReg_5_7,storeAddrNotKnownFlagsPReg_5_6,storeAddrNotKnownFlagsPReg_5_5,storeAddrNotKnownFlagsPReg_5_4,storeAddrNotKnownFlagsPReg_5_3,storeAddrNotKnownFlagsPReg_5_2,storeAddrNotKnownFlagsPReg_5_1,storeAddrNotKnownFlagsPReg_5_0}; // @[LoadQueue.scala 238:58:@9903.8]
  assign _T_25086 = {lastConflict_5_7,lastConflict_5_6,lastConflict_5_5,lastConflict_5_4,lastConflict_5_3,lastConflict_5_2,lastConflict_5_1,lastConflict_5_0}; // @[LoadQueue.scala 238:96:@9910.8]
  assign _T_25087 = _T_25079 < _T_25086; // @[LoadQueue.scala 238:61:@9911.8]
  assign _T_25088 = canBypass_5 & _T_25087; // @[LoadQueue.scala 237:64:@9912.8]
  assign _GEN_557 = _T_25049 ? _T_25088 : 1'h0; // @[LoadQueue.scala 230:110:@9876.6]
  assign bypassRequest_5 = _T_25041 ? _GEN_557 : 1'h0; // @[LoadQueue.scala 229:71:@9870.4]
  assign _GEN_530 = bypassRequest_5 ? 1'h1 : bypassInitiated_5; // @[LoadQueue.scala 217:34:@9599.6]
  assign _GEN_531 = initBits_5 ? 1'h0 : _GEN_530; // @[LoadQueue.scala 215:23:@9595.4]
  assign _T_25131 = {storeAddrNotKnownFlagsPReg_6_7,storeAddrNotKnownFlagsPReg_6_6,storeAddrNotKnownFlagsPReg_6_5,storeAddrNotKnownFlagsPReg_6_4,storeAddrNotKnownFlagsPReg_6_3,storeAddrNotKnownFlagsPReg_6_2,storeAddrNotKnownFlagsPReg_6_1,storeAddrNotKnownFlagsPReg_6_0}; // @[LoadQueue.scala 238:58:@9953.8]
  assign _T_25138 = {lastConflict_6_7,lastConflict_6_6,lastConflict_6_5,lastConflict_6_4,lastConflict_6_3,lastConflict_6_2,lastConflict_6_1,lastConflict_6_0}; // @[LoadQueue.scala 238:96:@9960.8]
  assign _T_25139 = _T_25131 < _T_25138; // @[LoadQueue.scala 238:61:@9961.8]
  assign _T_25140 = canBypass_6 & _T_25139; // @[LoadQueue.scala 237:64:@9962.8]
  assign _GEN_561 = _T_25101 ? _T_25140 : 1'h0; // @[LoadQueue.scala 230:110:@9926.6]
  assign bypassRequest_6 = _T_25093 ? _GEN_561 : 1'h0; // @[LoadQueue.scala 229:71:@9920.4]
  assign _GEN_532 = bypassRequest_6 ? 1'h1 : bypassInitiated_6; // @[LoadQueue.scala 217:34:@9606.6]
  assign _GEN_533 = initBits_6 ? 1'h0 : _GEN_532; // @[LoadQueue.scala 215:23:@9602.4]
  assign _T_25183 = {storeAddrNotKnownFlagsPReg_7_7,storeAddrNotKnownFlagsPReg_7_6,storeAddrNotKnownFlagsPReg_7_5,storeAddrNotKnownFlagsPReg_7_4,storeAddrNotKnownFlagsPReg_7_3,storeAddrNotKnownFlagsPReg_7_2,storeAddrNotKnownFlagsPReg_7_1,storeAddrNotKnownFlagsPReg_7_0}; // @[LoadQueue.scala 238:58:@10003.8]
  assign _T_25190 = {lastConflict_7_7,lastConflict_7_6,lastConflict_7_5,lastConflict_7_4,lastConflict_7_3,lastConflict_7_2,lastConflict_7_1,lastConflict_7_0}; // @[LoadQueue.scala 238:96:@10010.8]
  assign _T_25191 = _T_25183 < _T_25190; // @[LoadQueue.scala 238:61:@10011.8]
  assign _T_25192 = canBypass_7 & _T_25191; // @[LoadQueue.scala 237:64:@10012.8]
  assign _GEN_565 = _T_25153 ? _T_25192 : 1'h0; // @[LoadQueue.scala 230:110:@9976.6]
  assign bypassRequest_7 = _T_25145 ? _GEN_565 : 1'h0; // @[LoadQueue.scala 229:71:@9970.4]
  assign _GEN_534 = bypassRequest_7 ? 1'h1 : bypassInitiated_7; // @[LoadQueue.scala 217:34:@9613.6]
  assign _GEN_535 = initBits_7 ? 1'h0 : _GEN_534; // @[LoadQueue.scala 215:23:@9609.4]
  assign _T_25196 = loadRequest_0 | loadRequest_1; // @[LoadQueue.scala 247:28:@10018.4]
  assign _T_25197 = _T_25196 | loadRequest_2; // @[LoadQueue.scala 247:28:@10019.4]
  assign _T_25198 = _T_25197 | loadRequest_3; // @[LoadQueue.scala 247:28:@10020.4]
  assign _T_25199 = _T_25198 | loadRequest_4; // @[LoadQueue.scala 247:28:@10021.4]
  assign _T_25200 = _T_25199 | loadRequest_5; // @[LoadQueue.scala 247:28:@10022.4]
  assign _T_25201 = _T_25200 | loadRequest_6; // @[LoadQueue.scala 247:28:@10023.4]
  assign _T_25202 = _T_25201 | loadRequest_7; // @[LoadQueue.scala 247:28:@10024.4]
  assign _T_25211 = priorityLoadRequest_6 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@10026.6]
  assign _T_25212 = priorityLoadRequest_5 ? 3'h5 : _T_25211; // @[Mux.scala 31:69:@10027.6]
  assign _T_25213 = priorityLoadRequest_4 ? 3'h4 : _T_25212; // @[Mux.scala 31:69:@10028.6]
  assign _T_25214 = priorityLoadRequest_3 ? 3'h3 : _T_25213; // @[Mux.scala 31:69:@10029.6]
  assign _T_25215 = priorityLoadRequest_2 ? 3'h2 : _T_25214; // @[Mux.scala 31:69:@10030.6]
  assign _T_25216 = priorityLoadRequest_1 ? 3'h1 : _T_25215; // @[Mux.scala 31:69:@10031.6]
  assign _T_25217 = priorityLoadRequest_0 ? 3'h0 : _T_25216; // @[Mux.scala 31:69:@10032.6]
  assign _GEN_569 = 3'h1 == _T_25217 ? addrQ_1 : addrQ_0; // @[LoadQueue.scala 248:24:@10033.6]
  assign _GEN_570 = 3'h2 == _T_25217 ? addrQ_2 : _GEN_569; // @[LoadQueue.scala 248:24:@10033.6]
  assign _GEN_571 = 3'h3 == _T_25217 ? addrQ_3 : _GEN_570; // @[LoadQueue.scala 248:24:@10033.6]
  assign _GEN_572 = 3'h4 == _T_25217 ? addrQ_4 : _GEN_571; // @[LoadQueue.scala 248:24:@10033.6]
  assign _GEN_573 = 3'h5 == _T_25217 ? addrQ_5 : _GEN_572; // @[LoadQueue.scala 248:24:@10033.6]
  assign _GEN_574 = 3'h6 == _T_25217 ? addrQ_6 : _GEN_573; // @[LoadQueue.scala 248:24:@10033.6]
  assign _GEN_575 = 3'h7 == _T_25217 ? addrQ_7 : _GEN_574; // @[LoadQueue.scala 248:24:@10033.6]
  assign _T_25225 = prevPriorityRequest_0 | bypassRequest_0; // @[LoadQueue.scala 261:41:@10044.6]
  assign _GEN_578 = _T_25225 ? 1'h1 : dataKnown_0; // @[LoadQueue.scala 261:62:@10045.6]
  assign _GEN_579 = initBits_0 ? 1'h0 : _GEN_578; // @[LoadQueue.scala 259:25:@10040.4]
  assign _T_25228 = prevPriorityRequest_1 | bypassRequest_1; // @[LoadQueue.scala 261:41:@10052.6]
  assign _GEN_580 = _T_25228 ? 1'h1 : dataKnown_1; // @[LoadQueue.scala 261:62:@10053.6]
  assign _GEN_581 = initBits_1 ? 1'h0 : _GEN_580; // @[LoadQueue.scala 259:25:@10048.4]
  assign _T_25231 = prevPriorityRequest_2 | bypassRequest_2; // @[LoadQueue.scala 261:41:@10060.6]
  assign _GEN_582 = _T_25231 ? 1'h1 : dataKnown_2; // @[LoadQueue.scala 261:62:@10061.6]
  assign _GEN_583 = initBits_2 ? 1'h0 : _GEN_582; // @[LoadQueue.scala 259:25:@10056.4]
  assign _T_25234 = prevPriorityRequest_3 | bypassRequest_3; // @[LoadQueue.scala 261:41:@10068.6]
  assign _GEN_584 = _T_25234 ? 1'h1 : dataKnown_3; // @[LoadQueue.scala 261:62:@10069.6]
  assign _GEN_585 = initBits_3 ? 1'h0 : _GEN_584; // @[LoadQueue.scala 259:25:@10064.4]
  assign _T_25237 = prevPriorityRequest_4 | bypassRequest_4; // @[LoadQueue.scala 261:41:@10076.6]
  assign _GEN_586 = _T_25237 ? 1'h1 : dataKnown_4; // @[LoadQueue.scala 261:62:@10077.6]
  assign _GEN_587 = initBits_4 ? 1'h0 : _GEN_586; // @[LoadQueue.scala 259:25:@10072.4]
  assign _T_25240 = prevPriorityRequest_5 | bypassRequest_5; // @[LoadQueue.scala 261:41:@10084.6]
  assign _GEN_588 = _T_25240 ? 1'h1 : dataKnown_5; // @[LoadQueue.scala 261:62:@10085.6]
  assign _GEN_589 = initBits_5 ? 1'h0 : _GEN_588; // @[LoadQueue.scala 259:25:@10080.4]
  assign _T_25243 = prevPriorityRequest_6 | bypassRequest_6; // @[LoadQueue.scala 261:41:@10092.6]
  assign _GEN_590 = _T_25243 ? 1'h1 : dataKnown_6; // @[LoadQueue.scala 261:62:@10093.6]
  assign _GEN_591 = initBits_6 ? 1'h0 : _GEN_590; // @[LoadQueue.scala 259:25:@10088.4]
  assign _T_25246 = prevPriorityRequest_7 | bypassRequest_7; // @[LoadQueue.scala 261:41:@10100.6]
  assign _GEN_592 = _T_25246 ? 1'h1 : dataKnown_7; // @[LoadQueue.scala 261:62:@10101.6]
  assign _GEN_593 = initBits_7 ? 1'h0 : _GEN_592; // @[LoadQueue.scala 259:25:@10096.4]
  assign _GEN_594 = prevPriorityRequest_0 ? io_loadDataFromMem : dataQ_0; // @[LoadQueue.scala 269:44:@10108.6]
  assign _GEN_595 = bypassRequest_0 ? bypassVal_0 : _GEN_594; // @[LoadQueue.scala 267:32:@10104.4]
  assign _GEN_596 = prevPriorityRequest_1 ? io_loadDataFromMem : dataQ_1; // @[LoadQueue.scala 269:44:@10115.6]
  assign _GEN_597 = bypassRequest_1 ? bypassVal_1 : _GEN_596; // @[LoadQueue.scala 267:32:@10111.4]
  assign _GEN_598 = prevPriorityRequest_2 ? io_loadDataFromMem : dataQ_2; // @[LoadQueue.scala 269:44:@10122.6]
  assign _GEN_599 = bypassRequest_2 ? bypassVal_2 : _GEN_598; // @[LoadQueue.scala 267:32:@10118.4]
  assign _GEN_600 = prevPriorityRequest_3 ? io_loadDataFromMem : dataQ_3; // @[LoadQueue.scala 269:44:@10129.6]
  assign _GEN_601 = bypassRequest_3 ? bypassVal_3 : _GEN_600; // @[LoadQueue.scala 267:32:@10125.4]
  assign _GEN_602 = prevPriorityRequest_4 ? io_loadDataFromMem : dataQ_4; // @[LoadQueue.scala 269:44:@10136.6]
  assign _GEN_603 = bypassRequest_4 ? bypassVal_4 : _GEN_602; // @[LoadQueue.scala 267:32:@10132.4]
  assign _GEN_604 = prevPriorityRequest_5 ? io_loadDataFromMem : dataQ_5; // @[LoadQueue.scala 269:44:@10143.6]
  assign _GEN_605 = bypassRequest_5 ? bypassVal_5 : _GEN_604; // @[LoadQueue.scala 267:32:@10139.4]
  assign _GEN_606 = prevPriorityRequest_6 ? io_loadDataFromMem : dataQ_6; // @[LoadQueue.scala 269:44:@10150.6]
  assign _GEN_607 = bypassRequest_6 ? bypassVal_6 : _GEN_606; // @[LoadQueue.scala 267:32:@10146.4]
  assign _GEN_608 = prevPriorityRequest_7 ? io_loadDataFromMem : dataQ_7; // @[LoadQueue.scala 269:44:@10157.6]
  assign _GEN_609 = bypassRequest_7 ? bypassVal_7 : _GEN_608; // @[LoadQueue.scala 267:32:@10153.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[LoadQueue.scala 286:69:@10161.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[LoadQueue.scala 286:69:@10163.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[LoadQueue.scala 286:69:@10165.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[LoadQueue.scala 286:69:@10167.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[LoadQueue.scala 286:69:@10169.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[LoadQueue.scala 286:69:@10171.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[LoadQueue.scala 286:69:@10173.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[LoadQueue.scala 286:69:@10175.4]
  assign _T_25659 = addrKnown_0 == 1'h0; // @[LoadQueue.scala 298:86:@10195.4]
  assign _T_25660 = entriesPorts_0_0 & _T_25659; // @[LoadQueue.scala 298:83:@10196.4]
  assign _T_25662 = addrKnown_1 == 1'h0; // @[LoadQueue.scala 298:86:@10197.4]
  assign _T_25663 = entriesPorts_0_1 & _T_25662; // @[LoadQueue.scala 298:83:@10198.4]
  assign _T_25665 = addrKnown_2 == 1'h0; // @[LoadQueue.scala 298:86:@10199.4]
  assign _T_25666 = entriesPorts_0_2 & _T_25665; // @[LoadQueue.scala 298:83:@10200.4]
  assign _T_25668 = addrKnown_3 == 1'h0; // @[LoadQueue.scala 298:86:@10201.4]
  assign _T_25669 = entriesPorts_0_3 & _T_25668; // @[LoadQueue.scala 298:83:@10202.4]
  assign _T_25671 = addrKnown_4 == 1'h0; // @[LoadQueue.scala 298:86:@10203.4]
  assign _T_25672 = entriesPorts_0_4 & _T_25671; // @[LoadQueue.scala 298:83:@10204.4]
  assign _T_25674 = addrKnown_5 == 1'h0; // @[LoadQueue.scala 298:86:@10205.4]
  assign _T_25675 = entriesPorts_0_5 & _T_25674; // @[LoadQueue.scala 298:83:@10206.4]
  assign _T_25677 = addrKnown_6 == 1'h0; // @[LoadQueue.scala 298:86:@10207.4]
  assign _T_25678 = entriesPorts_0_6 & _T_25677; // @[LoadQueue.scala 298:83:@10208.4]
  assign _T_25680 = addrKnown_7 == 1'h0; // @[LoadQueue.scala 298:86:@10209.4]
  assign _T_25681 = entriesPorts_0_7 & _T_25680; // @[LoadQueue.scala 298:83:@10210.4]
  assign _T_25732 = _T_25681 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10240.4]
  assign _T_25733 = _T_25678 ? 8'h40 : _T_25732; // @[Mux.scala 31:69:@10241.4]
  assign _T_25734 = _T_25675 ? 8'h20 : _T_25733; // @[Mux.scala 31:69:@10242.4]
  assign _T_25735 = _T_25672 ? 8'h10 : _T_25734; // @[Mux.scala 31:69:@10243.4]
  assign _T_25736 = _T_25669 ? 8'h8 : _T_25735; // @[Mux.scala 31:69:@10244.4]
  assign _T_25737 = _T_25666 ? 8'h4 : _T_25736; // @[Mux.scala 31:69:@10245.4]
  assign _T_25738 = _T_25663 ? 8'h2 : _T_25737; // @[Mux.scala 31:69:@10246.4]
  assign _T_25739 = _T_25660 ? 8'h1 : _T_25738; // @[Mux.scala 31:69:@10247.4]
  assign _T_25740 = _T_25739[0]; // @[OneHot.scala 66:30:@10248.4]
  assign _T_25741 = _T_25739[1]; // @[OneHot.scala 66:30:@10249.4]
  assign _T_25742 = _T_25739[2]; // @[OneHot.scala 66:30:@10250.4]
  assign _T_25743 = _T_25739[3]; // @[OneHot.scala 66:30:@10251.4]
  assign _T_25744 = _T_25739[4]; // @[OneHot.scala 66:30:@10252.4]
  assign _T_25745 = _T_25739[5]; // @[OneHot.scala 66:30:@10253.4]
  assign _T_25746 = _T_25739[6]; // @[OneHot.scala 66:30:@10254.4]
  assign _T_25747 = _T_25739[7]; // @[OneHot.scala 66:30:@10255.4]
  assign _T_25772 = _T_25660 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10265.4]
  assign _T_25773 = _T_25681 ? 8'h40 : _T_25772; // @[Mux.scala 31:69:@10266.4]
  assign _T_25774 = _T_25678 ? 8'h20 : _T_25773; // @[Mux.scala 31:69:@10267.4]
  assign _T_25775 = _T_25675 ? 8'h10 : _T_25774; // @[Mux.scala 31:69:@10268.4]
  assign _T_25776 = _T_25672 ? 8'h8 : _T_25775; // @[Mux.scala 31:69:@10269.4]
  assign _T_25777 = _T_25669 ? 8'h4 : _T_25776; // @[Mux.scala 31:69:@10270.4]
  assign _T_25778 = _T_25666 ? 8'h2 : _T_25777; // @[Mux.scala 31:69:@10271.4]
  assign _T_25779 = _T_25663 ? 8'h1 : _T_25778; // @[Mux.scala 31:69:@10272.4]
  assign _T_25780 = _T_25779[0]; // @[OneHot.scala 66:30:@10273.4]
  assign _T_25781 = _T_25779[1]; // @[OneHot.scala 66:30:@10274.4]
  assign _T_25782 = _T_25779[2]; // @[OneHot.scala 66:30:@10275.4]
  assign _T_25783 = _T_25779[3]; // @[OneHot.scala 66:30:@10276.4]
  assign _T_25784 = _T_25779[4]; // @[OneHot.scala 66:30:@10277.4]
  assign _T_25785 = _T_25779[5]; // @[OneHot.scala 66:30:@10278.4]
  assign _T_25786 = _T_25779[6]; // @[OneHot.scala 66:30:@10279.4]
  assign _T_25787 = _T_25779[7]; // @[OneHot.scala 66:30:@10280.4]
  assign _T_25812 = _T_25663 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10290.4]
  assign _T_25813 = _T_25660 ? 8'h40 : _T_25812; // @[Mux.scala 31:69:@10291.4]
  assign _T_25814 = _T_25681 ? 8'h20 : _T_25813; // @[Mux.scala 31:69:@10292.4]
  assign _T_25815 = _T_25678 ? 8'h10 : _T_25814; // @[Mux.scala 31:69:@10293.4]
  assign _T_25816 = _T_25675 ? 8'h8 : _T_25815; // @[Mux.scala 31:69:@10294.4]
  assign _T_25817 = _T_25672 ? 8'h4 : _T_25816; // @[Mux.scala 31:69:@10295.4]
  assign _T_25818 = _T_25669 ? 8'h2 : _T_25817; // @[Mux.scala 31:69:@10296.4]
  assign _T_25819 = _T_25666 ? 8'h1 : _T_25818; // @[Mux.scala 31:69:@10297.4]
  assign _T_25820 = _T_25819[0]; // @[OneHot.scala 66:30:@10298.4]
  assign _T_25821 = _T_25819[1]; // @[OneHot.scala 66:30:@10299.4]
  assign _T_25822 = _T_25819[2]; // @[OneHot.scala 66:30:@10300.4]
  assign _T_25823 = _T_25819[3]; // @[OneHot.scala 66:30:@10301.4]
  assign _T_25824 = _T_25819[4]; // @[OneHot.scala 66:30:@10302.4]
  assign _T_25825 = _T_25819[5]; // @[OneHot.scala 66:30:@10303.4]
  assign _T_25826 = _T_25819[6]; // @[OneHot.scala 66:30:@10304.4]
  assign _T_25827 = _T_25819[7]; // @[OneHot.scala 66:30:@10305.4]
  assign _T_25852 = _T_25666 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10315.4]
  assign _T_25853 = _T_25663 ? 8'h40 : _T_25852; // @[Mux.scala 31:69:@10316.4]
  assign _T_25854 = _T_25660 ? 8'h20 : _T_25853; // @[Mux.scala 31:69:@10317.4]
  assign _T_25855 = _T_25681 ? 8'h10 : _T_25854; // @[Mux.scala 31:69:@10318.4]
  assign _T_25856 = _T_25678 ? 8'h8 : _T_25855; // @[Mux.scala 31:69:@10319.4]
  assign _T_25857 = _T_25675 ? 8'h4 : _T_25856; // @[Mux.scala 31:69:@10320.4]
  assign _T_25858 = _T_25672 ? 8'h2 : _T_25857; // @[Mux.scala 31:69:@10321.4]
  assign _T_25859 = _T_25669 ? 8'h1 : _T_25858; // @[Mux.scala 31:69:@10322.4]
  assign _T_25860 = _T_25859[0]; // @[OneHot.scala 66:30:@10323.4]
  assign _T_25861 = _T_25859[1]; // @[OneHot.scala 66:30:@10324.4]
  assign _T_25862 = _T_25859[2]; // @[OneHot.scala 66:30:@10325.4]
  assign _T_25863 = _T_25859[3]; // @[OneHot.scala 66:30:@10326.4]
  assign _T_25864 = _T_25859[4]; // @[OneHot.scala 66:30:@10327.4]
  assign _T_25865 = _T_25859[5]; // @[OneHot.scala 66:30:@10328.4]
  assign _T_25866 = _T_25859[6]; // @[OneHot.scala 66:30:@10329.4]
  assign _T_25867 = _T_25859[7]; // @[OneHot.scala 66:30:@10330.4]
  assign _T_25892 = _T_25669 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10340.4]
  assign _T_25893 = _T_25666 ? 8'h40 : _T_25892; // @[Mux.scala 31:69:@10341.4]
  assign _T_25894 = _T_25663 ? 8'h20 : _T_25893; // @[Mux.scala 31:69:@10342.4]
  assign _T_25895 = _T_25660 ? 8'h10 : _T_25894; // @[Mux.scala 31:69:@10343.4]
  assign _T_25896 = _T_25681 ? 8'h8 : _T_25895; // @[Mux.scala 31:69:@10344.4]
  assign _T_25897 = _T_25678 ? 8'h4 : _T_25896; // @[Mux.scala 31:69:@10345.4]
  assign _T_25898 = _T_25675 ? 8'h2 : _T_25897; // @[Mux.scala 31:69:@10346.4]
  assign _T_25899 = _T_25672 ? 8'h1 : _T_25898; // @[Mux.scala 31:69:@10347.4]
  assign _T_25900 = _T_25899[0]; // @[OneHot.scala 66:30:@10348.4]
  assign _T_25901 = _T_25899[1]; // @[OneHot.scala 66:30:@10349.4]
  assign _T_25902 = _T_25899[2]; // @[OneHot.scala 66:30:@10350.4]
  assign _T_25903 = _T_25899[3]; // @[OneHot.scala 66:30:@10351.4]
  assign _T_25904 = _T_25899[4]; // @[OneHot.scala 66:30:@10352.4]
  assign _T_25905 = _T_25899[5]; // @[OneHot.scala 66:30:@10353.4]
  assign _T_25906 = _T_25899[6]; // @[OneHot.scala 66:30:@10354.4]
  assign _T_25907 = _T_25899[7]; // @[OneHot.scala 66:30:@10355.4]
  assign _T_25932 = _T_25672 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10365.4]
  assign _T_25933 = _T_25669 ? 8'h40 : _T_25932; // @[Mux.scala 31:69:@10366.4]
  assign _T_25934 = _T_25666 ? 8'h20 : _T_25933; // @[Mux.scala 31:69:@10367.4]
  assign _T_25935 = _T_25663 ? 8'h10 : _T_25934; // @[Mux.scala 31:69:@10368.4]
  assign _T_25936 = _T_25660 ? 8'h8 : _T_25935; // @[Mux.scala 31:69:@10369.4]
  assign _T_25937 = _T_25681 ? 8'h4 : _T_25936; // @[Mux.scala 31:69:@10370.4]
  assign _T_25938 = _T_25678 ? 8'h2 : _T_25937; // @[Mux.scala 31:69:@10371.4]
  assign _T_25939 = _T_25675 ? 8'h1 : _T_25938; // @[Mux.scala 31:69:@10372.4]
  assign _T_25940 = _T_25939[0]; // @[OneHot.scala 66:30:@10373.4]
  assign _T_25941 = _T_25939[1]; // @[OneHot.scala 66:30:@10374.4]
  assign _T_25942 = _T_25939[2]; // @[OneHot.scala 66:30:@10375.4]
  assign _T_25943 = _T_25939[3]; // @[OneHot.scala 66:30:@10376.4]
  assign _T_25944 = _T_25939[4]; // @[OneHot.scala 66:30:@10377.4]
  assign _T_25945 = _T_25939[5]; // @[OneHot.scala 66:30:@10378.4]
  assign _T_25946 = _T_25939[6]; // @[OneHot.scala 66:30:@10379.4]
  assign _T_25947 = _T_25939[7]; // @[OneHot.scala 66:30:@10380.4]
  assign _T_25972 = _T_25675 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10390.4]
  assign _T_25973 = _T_25672 ? 8'h40 : _T_25972; // @[Mux.scala 31:69:@10391.4]
  assign _T_25974 = _T_25669 ? 8'h20 : _T_25973; // @[Mux.scala 31:69:@10392.4]
  assign _T_25975 = _T_25666 ? 8'h10 : _T_25974; // @[Mux.scala 31:69:@10393.4]
  assign _T_25976 = _T_25663 ? 8'h8 : _T_25975; // @[Mux.scala 31:69:@10394.4]
  assign _T_25977 = _T_25660 ? 8'h4 : _T_25976; // @[Mux.scala 31:69:@10395.4]
  assign _T_25978 = _T_25681 ? 8'h2 : _T_25977; // @[Mux.scala 31:69:@10396.4]
  assign _T_25979 = _T_25678 ? 8'h1 : _T_25978; // @[Mux.scala 31:69:@10397.4]
  assign _T_25980 = _T_25979[0]; // @[OneHot.scala 66:30:@10398.4]
  assign _T_25981 = _T_25979[1]; // @[OneHot.scala 66:30:@10399.4]
  assign _T_25982 = _T_25979[2]; // @[OneHot.scala 66:30:@10400.4]
  assign _T_25983 = _T_25979[3]; // @[OneHot.scala 66:30:@10401.4]
  assign _T_25984 = _T_25979[4]; // @[OneHot.scala 66:30:@10402.4]
  assign _T_25985 = _T_25979[5]; // @[OneHot.scala 66:30:@10403.4]
  assign _T_25986 = _T_25979[6]; // @[OneHot.scala 66:30:@10404.4]
  assign _T_25987 = _T_25979[7]; // @[OneHot.scala 66:30:@10405.4]
  assign _T_26012 = _T_25678 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10415.4]
  assign _T_26013 = _T_25675 ? 8'h40 : _T_26012; // @[Mux.scala 31:69:@10416.4]
  assign _T_26014 = _T_25672 ? 8'h20 : _T_26013; // @[Mux.scala 31:69:@10417.4]
  assign _T_26015 = _T_25669 ? 8'h10 : _T_26014; // @[Mux.scala 31:69:@10418.4]
  assign _T_26016 = _T_25666 ? 8'h8 : _T_26015; // @[Mux.scala 31:69:@10419.4]
  assign _T_26017 = _T_25663 ? 8'h4 : _T_26016; // @[Mux.scala 31:69:@10420.4]
  assign _T_26018 = _T_25660 ? 8'h2 : _T_26017; // @[Mux.scala 31:69:@10421.4]
  assign _T_26019 = _T_25681 ? 8'h1 : _T_26018; // @[Mux.scala 31:69:@10422.4]
  assign _T_26020 = _T_26019[0]; // @[OneHot.scala 66:30:@10423.4]
  assign _T_26021 = _T_26019[1]; // @[OneHot.scala 66:30:@10424.4]
  assign _T_26022 = _T_26019[2]; // @[OneHot.scala 66:30:@10425.4]
  assign _T_26023 = _T_26019[3]; // @[OneHot.scala 66:30:@10426.4]
  assign _T_26024 = _T_26019[4]; // @[OneHot.scala 66:30:@10427.4]
  assign _T_26025 = _T_26019[5]; // @[OneHot.scala 66:30:@10428.4]
  assign _T_26026 = _T_26019[6]; // @[OneHot.scala 66:30:@10429.4]
  assign _T_26027 = _T_26019[7]; // @[OneHot.scala 66:30:@10430.4]
  assign _T_26068 = {_T_25747,_T_25746,_T_25745,_T_25744,_T_25743,_T_25742,_T_25741,_T_25740}; // @[Mux.scala 19:72:@10446.4]
  assign _T_26070 = _T_24152 ? _T_26068 : 8'h0; // @[Mux.scala 19:72:@10447.4]
  assign _T_26077 = {_T_25786,_T_25785,_T_25784,_T_25783,_T_25782,_T_25781,_T_25780,_T_25787}; // @[Mux.scala 19:72:@10454.4]
  assign _T_26079 = _T_24153 ? _T_26077 : 8'h0; // @[Mux.scala 19:72:@10455.4]
  assign _T_26086 = {_T_25825,_T_25824,_T_25823,_T_25822,_T_25821,_T_25820,_T_25827,_T_25826}; // @[Mux.scala 19:72:@10462.4]
  assign _T_26088 = _T_24154 ? _T_26086 : 8'h0; // @[Mux.scala 19:72:@10463.4]
  assign _T_26095 = {_T_25864,_T_25863,_T_25862,_T_25861,_T_25860,_T_25867,_T_25866,_T_25865}; // @[Mux.scala 19:72:@10470.4]
  assign _T_26097 = _T_24155 ? _T_26095 : 8'h0; // @[Mux.scala 19:72:@10471.4]
  assign _T_26104 = {_T_25903,_T_25902,_T_25901,_T_25900,_T_25907,_T_25906,_T_25905,_T_25904}; // @[Mux.scala 19:72:@10478.4]
  assign _T_26106 = _T_24156 ? _T_26104 : 8'h0; // @[Mux.scala 19:72:@10479.4]
  assign _T_26113 = {_T_25942,_T_25941,_T_25940,_T_25947,_T_25946,_T_25945,_T_25944,_T_25943}; // @[Mux.scala 19:72:@10486.4]
  assign _T_26115 = _T_24157 ? _T_26113 : 8'h0; // @[Mux.scala 19:72:@10487.4]
  assign _T_26122 = {_T_25981,_T_25980,_T_25987,_T_25986,_T_25985,_T_25984,_T_25983,_T_25982}; // @[Mux.scala 19:72:@10494.4]
  assign _T_26124 = _T_24158 ? _T_26122 : 8'h0; // @[Mux.scala 19:72:@10495.4]
  assign _T_26131 = {_T_26020,_T_26027,_T_26026,_T_26025,_T_26024,_T_26023,_T_26022,_T_26021}; // @[Mux.scala 19:72:@10502.4]
  assign _T_26133 = _T_24159 ? _T_26131 : 8'h0; // @[Mux.scala 19:72:@10503.4]
  assign _T_26134 = _T_26070 | _T_26079; // @[Mux.scala 19:72:@10504.4]
  assign _T_26135 = _T_26134 | _T_26088; // @[Mux.scala 19:72:@10505.4]
  assign _T_26136 = _T_26135 | _T_26097; // @[Mux.scala 19:72:@10506.4]
  assign _T_26137 = _T_26136 | _T_26106; // @[Mux.scala 19:72:@10507.4]
  assign _T_26138 = _T_26137 | _T_26115; // @[Mux.scala 19:72:@10508.4]
  assign _T_26139 = _T_26138 | _T_26124; // @[Mux.scala 19:72:@10509.4]
  assign _T_26140 = _T_26139 | _T_26133; // @[Mux.scala 19:72:@10510.4]
  assign inputPriorityPorts_0_0 = _T_26140[0]; // @[Mux.scala 19:72:@10514.4]
  assign inputPriorityPorts_0_1 = _T_26140[1]; // @[Mux.scala 19:72:@10516.4]
  assign inputPriorityPorts_0_2 = _T_26140[2]; // @[Mux.scala 19:72:@10518.4]
  assign inputPriorityPorts_0_3 = _T_26140[3]; // @[Mux.scala 19:72:@10520.4]
  assign inputPriorityPorts_0_4 = _T_26140[4]; // @[Mux.scala 19:72:@10522.4]
  assign inputPriorityPorts_0_5 = _T_26140[5]; // @[Mux.scala 19:72:@10524.4]
  assign inputPriorityPorts_0_6 = _T_26140[6]; // @[Mux.scala 19:72:@10526.4]
  assign inputPriorityPorts_0_7 = _T_26140[7]; // @[Mux.scala 19:72:@10528.4]
  assign _T_26254 = entriesPorts_0_7 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10558.4]
  assign _T_26255 = entriesPorts_0_6 ? 8'h40 : _T_26254; // @[Mux.scala 31:69:@10559.4]
  assign _T_26256 = entriesPorts_0_5 ? 8'h20 : _T_26255; // @[Mux.scala 31:69:@10560.4]
  assign _T_26257 = entriesPorts_0_4 ? 8'h10 : _T_26256; // @[Mux.scala 31:69:@10561.4]
  assign _T_26258 = entriesPorts_0_3 ? 8'h8 : _T_26257; // @[Mux.scala 31:69:@10562.4]
  assign _T_26259 = entriesPorts_0_2 ? 8'h4 : _T_26258; // @[Mux.scala 31:69:@10563.4]
  assign _T_26260 = entriesPorts_0_1 ? 8'h2 : _T_26259; // @[Mux.scala 31:69:@10564.4]
  assign _T_26261 = entriesPorts_0_0 ? 8'h1 : _T_26260; // @[Mux.scala 31:69:@10565.4]
  assign _T_26262 = _T_26261[0]; // @[OneHot.scala 66:30:@10566.4]
  assign _T_26263 = _T_26261[1]; // @[OneHot.scala 66:30:@10567.4]
  assign _T_26264 = _T_26261[2]; // @[OneHot.scala 66:30:@10568.4]
  assign _T_26265 = _T_26261[3]; // @[OneHot.scala 66:30:@10569.4]
  assign _T_26266 = _T_26261[4]; // @[OneHot.scala 66:30:@10570.4]
  assign _T_26267 = _T_26261[5]; // @[OneHot.scala 66:30:@10571.4]
  assign _T_26268 = _T_26261[6]; // @[OneHot.scala 66:30:@10572.4]
  assign _T_26269 = _T_26261[7]; // @[OneHot.scala 66:30:@10573.4]
  assign _T_26294 = entriesPorts_0_0 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10583.4]
  assign _T_26295 = entriesPorts_0_7 ? 8'h40 : _T_26294; // @[Mux.scala 31:69:@10584.4]
  assign _T_26296 = entriesPorts_0_6 ? 8'h20 : _T_26295; // @[Mux.scala 31:69:@10585.4]
  assign _T_26297 = entriesPorts_0_5 ? 8'h10 : _T_26296; // @[Mux.scala 31:69:@10586.4]
  assign _T_26298 = entriesPorts_0_4 ? 8'h8 : _T_26297; // @[Mux.scala 31:69:@10587.4]
  assign _T_26299 = entriesPorts_0_3 ? 8'h4 : _T_26298; // @[Mux.scala 31:69:@10588.4]
  assign _T_26300 = entriesPorts_0_2 ? 8'h2 : _T_26299; // @[Mux.scala 31:69:@10589.4]
  assign _T_26301 = entriesPorts_0_1 ? 8'h1 : _T_26300; // @[Mux.scala 31:69:@10590.4]
  assign _T_26302 = _T_26301[0]; // @[OneHot.scala 66:30:@10591.4]
  assign _T_26303 = _T_26301[1]; // @[OneHot.scala 66:30:@10592.4]
  assign _T_26304 = _T_26301[2]; // @[OneHot.scala 66:30:@10593.4]
  assign _T_26305 = _T_26301[3]; // @[OneHot.scala 66:30:@10594.4]
  assign _T_26306 = _T_26301[4]; // @[OneHot.scala 66:30:@10595.4]
  assign _T_26307 = _T_26301[5]; // @[OneHot.scala 66:30:@10596.4]
  assign _T_26308 = _T_26301[6]; // @[OneHot.scala 66:30:@10597.4]
  assign _T_26309 = _T_26301[7]; // @[OneHot.scala 66:30:@10598.4]
  assign _T_26334 = entriesPorts_0_1 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10608.4]
  assign _T_26335 = entriesPorts_0_0 ? 8'h40 : _T_26334; // @[Mux.scala 31:69:@10609.4]
  assign _T_26336 = entriesPorts_0_7 ? 8'h20 : _T_26335; // @[Mux.scala 31:69:@10610.4]
  assign _T_26337 = entriesPorts_0_6 ? 8'h10 : _T_26336; // @[Mux.scala 31:69:@10611.4]
  assign _T_26338 = entriesPorts_0_5 ? 8'h8 : _T_26337; // @[Mux.scala 31:69:@10612.4]
  assign _T_26339 = entriesPorts_0_4 ? 8'h4 : _T_26338; // @[Mux.scala 31:69:@10613.4]
  assign _T_26340 = entriesPorts_0_3 ? 8'h2 : _T_26339; // @[Mux.scala 31:69:@10614.4]
  assign _T_26341 = entriesPorts_0_2 ? 8'h1 : _T_26340; // @[Mux.scala 31:69:@10615.4]
  assign _T_26342 = _T_26341[0]; // @[OneHot.scala 66:30:@10616.4]
  assign _T_26343 = _T_26341[1]; // @[OneHot.scala 66:30:@10617.4]
  assign _T_26344 = _T_26341[2]; // @[OneHot.scala 66:30:@10618.4]
  assign _T_26345 = _T_26341[3]; // @[OneHot.scala 66:30:@10619.4]
  assign _T_26346 = _T_26341[4]; // @[OneHot.scala 66:30:@10620.4]
  assign _T_26347 = _T_26341[5]; // @[OneHot.scala 66:30:@10621.4]
  assign _T_26348 = _T_26341[6]; // @[OneHot.scala 66:30:@10622.4]
  assign _T_26349 = _T_26341[7]; // @[OneHot.scala 66:30:@10623.4]
  assign _T_26374 = entriesPorts_0_2 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10633.4]
  assign _T_26375 = entriesPorts_0_1 ? 8'h40 : _T_26374; // @[Mux.scala 31:69:@10634.4]
  assign _T_26376 = entriesPorts_0_0 ? 8'h20 : _T_26375; // @[Mux.scala 31:69:@10635.4]
  assign _T_26377 = entriesPorts_0_7 ? 8'h10 : _T_26376; // @[Mux.scala 31:69:@10636.4]
  assign _T_26378 = entriesPorts_0_6 ? 8'h8 : _T_26377; // @[Mux.scala 31:69:@10637.4]
  assign _T_26379 = entriesPorts_0_5 ? 8'h4 : _T_26378; // @[Mux.scala 31:69:@10638.4]
  assign _T_26380 = entriesPorts_0_4 ? 8'h2 : _T_26379; // @[Mux.scala 31:69:@10639.4]
  assign _T_26381 = entriesPorts_0_3 ? 8'h1 : _T_26380; // @[Mux.scala 31:69:@10640.4]
  assign _T_26382 = _T_26381[0]; // @[OneHot.scala 66:30:@10641.4]
  assign _T_26383 = _T_26381[1]; // @[OneHot.scala 66:30:@10642.4]
  assign _T_26384 = _T_26381[2]; // @[OneHot.scala 66:30:@10643.4]
  assign _T_26385 = _T_26381[3]; // @[OneHot.scala 66:30:@10644.4]
  assign _T_26386 = _T_26381[4]; // @[OneHot.scala 66:30:@10645.4]
  assign _T_26387 = _T_26381[5]; // @[OneHot.scala 66:30:@10646.4]
  assign _T_26388 = _T_26381[6]; // @[OneHot.scala 66:30:@10647.4]
  assign _T_26389 = _T_26381[7]; // @[OneHot.scala 66:30:@10648.4]
  assign _T_26414 = entriesPorts_0_3 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10658.4]
  assign _T_26415 = entriesPorts_0_2 ? 8'h40 : _T_26414; // @[Mux.scala 31:69:@10659.4]
  assign _T_26416 = entriesPorts_0_1 ? 8'h20 : _T_26415; // @[Mux.scala 31:69:@10660.4]
  assign _T_26417 = entriesPorts_0_0 ? 8'h10 : _T_26416; // @[Mux.scala 31:69:@10661.4]
  assign _T_26418 = entriesPorts_0_7 ? 8'h8 : _T_26417; // @[Mux.scala 31:69:@10662.4]
  assign _T_26419 = entriesPorts_0_6 ? 8'h4 : _T_26418; // @[Mux.scala 31:69:@10663.4]
  assign _T_26420 = entriesPorts_0_5 ? 8'h2 : _T_26419; // @[Mux.scala 31:69:@10664.4]
  assign _T_26421 = entriesPorts_0_4 ? 8'h1 : _T_26420; // @[Mux.scala 31:69:@10665.4]
  assign _T_26422 = _T_26421[0]; // @[OneHot.scala 66:30:@10666.4]
  assign _T_26423 = _T_26421[1]; // @[OneHot.scala 66:30:@10667.4]
  assign _T_26424 = _T_26421[2]; // @[OneHot.scala 66:30:@10668.4]
  assign _T_26425 = _T_26421[3]; // @[OneHot.scala 66:30:@10669.4]
  assign _T_26426 = _T_26421[4]; // @[OneHot.scala 66:30:@10670.4]
  assign _T_26427 = _T_26421[5]; // @[OneHot.scala 66:30:@10671.4]
  assign _T_26428 = _T_26421[6]; // @[OneHot.scala 66:30:@10672.4]
  assign _T_26429 = _T_26421[7]; // @[OneHot.scala 66:30:@10673.4]
  assign _T_26454 = entriesPorts_0_4 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10683.4]
  assign _T_26455 = entriesPorts_0_3 ? 8'h40 : _T_26454; // @[Mux.scala 31:69:@10684.4]
  assign _T_26456 = entriesPorts_0_2 ? 8'h20 : _T_26455; // @[Mux.scala 31:69:@10685.4]
  assign _T_26457 = entriesPorts_0_1 ? 8'h10 : _T_26456; // @[Mux.scala 31:69:@10686.4]
  assign _T_26458 = entriesPorts_0_0 ? 8'h8 : _T_26457; // @[Mux.scala 31:69:@10687.4]
  assign _T_26459 = entriesPorts_0_7 ? 8'h4 : _T_26458; // @[Mux.scala 31:69:@10688.4]
  assign _T_26460 = entriesPorts_0_6 ? 8'h2 : _T_26459; // @[Mux.scala 31:69:@10689.4]
  assign _T_26461 = entriesPorts_0_5 ? 8'h1 : _T_26460; // @[Mux.scala 31:69:@10690.4]
  assign _T_26462 = _T_26461[0]; // @[OneHot.scala 66:30:@10691.4]
  assign _T_26463 = _T_26461[1]; // @[OneHot.scala 66:30:@10692.4]
  assign _T_26464 = _T_26461[2]; // @[OneHot.scala 66:30:@10693.4]
  assign _T_26465 = _T_26461[3]; // @[OneHot.scala 66:30:@10694.4]
  assign _T_26466 = _T_26461[4]; // @[OneHot.scala 66:30:@10695.4]
  assign _T_26467 = _T_26461[5]; // @[OneHot.scala 66:30:@10696.4]
  assign _T_26468 = _T_26461[6]; // @[OneHot.scala 66:30:@10697.4]
  assign _T_26469 = _T_26461[7]; // @[OneHot.scala 66:30:@10698.4]
  assign _T_26494 = entriesPorts_0_5 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10708.4]
  assign _T_26495 = entriesPorts_0_4 ? 8'h40 : _T_26494; // @[Mux.scala 31:69:@10709.4]
  assign _T_26496 = entriesPorts_0_3 ? 8'h20 : _T_26495; // @[Mux.scala 31:69:@10710.4]
  assign _T_26497 = entriesPorts_0_2 ? 8'h10 : _T_26496; // @[Mux.scala 31:69:@10711.4]
  assign _T_26498 = entriesPorts_0_1 ? 8'h8 : _T_26497; // @[Mux.scala 31:69:@10712.4]
  assign _T_26499 = entriesPorts_0_0 ? 8'h4 : _T_26498; // @[Mux.scala 31:69:@10713.4]
  assign _T_26500 = entriesPorts_0_7 ? 8'h2 : _T_26499; // @[Mux.scala 31:69:@10714.4]
  assign _T_26501 = entriesPorts_0_6 ? 8'h1 : _T_26500; // @[Mux.scala 31:69:@10715.4]
  assign _T_26502 = _T_26501[0]; // @[OneHot.scala 66:30:@10716.4]
  assign _T_26503 = _T_26501[1]; // @[OneHot.scala 66:30:@10717.4]
  assign _T_26504 = _T_26501[2]; // @[OneHot.scala 66:30:@10718.4]
  assign _T_26505 = _T_26501[3]; // @[OneHot.scala 66:30:@10719.4]
  assign _T_26506 = _T_26501[4]; // @[OneHot.scala 66:30:@10720.4]
  assign _T_26507 = _T_26501[5]; // @[OneHot.scala 66:30:@10721.4]
  assign _T_26508 = _T_26501[6]; // @[OneHot.scala 66:30:@10722.4]
  assign _T_26509 = _T_26501[7]; // @[OneHot.scala 66:30:@10723.4]
  assign _T_26534 = entriesPorts_0_6 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10733.4]
  assign _T_26535 = entriesPorts_0_5 ? 8'h40 : _T_26534; // @[Mux.scala 31:69:@10734.4]
  assign _T_26536 = entriesPorts_0_4 ? 8'h20 : _T_26535; // @[Mux.scala 31:69:@10735.4]
  assign _T_26537 = entriesPorts_0_3 ? 8'h10 : _T_26536; // @[Mux.scala 31:69:@10736.4]
  assign _T_26538 = entriesPorts_0_2 ? 8'h8 : _T_26537; // @[Mux.scala 31:69:@10737.4]
  assign _T_26539 = entriesPorts_0_1 ? 8'h4 : _T_26538; // @[Mux.scala 31:69:@10738.4]
  assign _T_26540 = entriesPorts_0_0 ? 8'h2 : _T_26539; // @[Mux.scala 31:69:@10739.4]
  assign _T_26541 = entriesPorts_0_7 ? 8'h1 : _T_26540; // @[Mux.scala 31:69:@10740.4]
  assign _T_26542 = _T_26541[0]; // @[OneHot.scala 66:30:@10741.4]
  assign _T_26543 = _T_26541[1]; // @[OneHot.scala 66:30:@10742.4]
  assign _T_26544 = _T_26541[2]; // @[OneHot.scala 66:30:@10743.4]
  assign _T_26545 = _T_26541[3]; // @[OneHot.scala 66:30:@10744.4]
  assign _T_26546 = _T_26541[4]; // @[OneHot.scala 66:30:@10745.4]
  assign _T_26547 = _T_26541[5]; // @[OneHot.scala 66:30:@10746.4]
  assign _T_26548 = _T_26541[6]; // @[OneHot.scala 66:30:@10747.4]
  assign _T_26549 = _T_26541[7]; // @[OneHot.scala 66:30:@10748.4]
  assign _T_26590 = {_T_26269,_T_26268,_T_26267,_T_26266,_T_26265,_T_26264,_T_26263,_T_26262}; // @[Mux.scala 19:72:@10764.4]
  assign _T_26592 = _T_24152 ? _T_26590 : 8'h0; // @[Mux.scala 19:72:@10765.4]
  assign _T_26599 = {_T_26308,_T_26307,_T_26306,_T_26305,_T_26304,_T_26303,_T_26302,_T_26309}; // @[Mux.scala 19:72:@10772.4]
  assign _T_26601 = _T_24153 ? _T_26599 : 8'h0; // @[Mux.scala 19:72:@10773.4]
  assign _T_26608 = {_T_26347,_T_26346,_T_26345,_T_26344,_T_26343,_T_26342,_T_26349,_T_26348}; // @[Mux.scala 19:72:@10780.4]
  assign _T_26610 = _T_24154 ? _T_26608 : 8'h0; // @[Mux.scala 19:72:@10781.4]
  assign _T_26617 = {_T_26386,_T_26385,_T_26384,_T_26383,_T_26382,_T_26389,_T_26388,_T_26387}; // @[Mux.scala 19:72:@10788.4]
  assign _T_26619 = _T_24155 ? _T_26617 : 8'h0; // @[Mux.scala 19:72:@10789.4]
  assign _T_26626 = {_T_26425,_T_26424,_T_26423,_T_26422,_T_26429,_T_26428,_T_26427,_T_26426}; // @[Mux.scala 19:72:@10796.4]
  assign _T_26628 = _T_24156 ? _T_26626 : 8'h0; // @[Mux.scala 19:72:@10797.4]
  assign _T_26635 = {_T_26464,_T_26463,_T_26462,_T_26469,_T_26468,_T_26467,_T_26466,_T_26465}; // @[Mux.scala 19:72:@10804.4]
  assign _T_26637 = _T_24157 ? _T_26635 : 8'h0; // @[Mux.scala 19:72:@10805.4]
  assign _T_26644 = {_T_26503,_T_26502,_T_26509,_T_26508,_T_26507,_T_26506,_T_26505,_T_26504}; // @[Mux.scala 19:72:@10812.4]
  assign _T_26646 = _T_24158 ? _T_26644 : 8'h0; // @[Mux.scala 19:72:@10813.4]
  assign _T_26653 = {_T_26542,_T_26549,_T_26548,_T_26547,_T_26546,_T_26545,_T_26544,_T_26543}; // @[Mux.scala 19:72:@10820.4]
  assign _T_26655 = _T_24159 ? _T_26653 : 8'h0; // @[Mux.scala 19:72:@10821.4]
  assign _T_26656 = _T_26592 | _T_26601; // @[Mux.scala 19:72:@10822.4]
  assign _T_26657 = _T_26656 | _T_26610; // @[Mux.scala 19:72:@10823.4]
  assign _T_26658 = _T_26657 | _T_26619; // @[Mux.scala 19:72:@10824.4]
  assign _T_26659 = _T_26658 | _T_26628; // @[Mux.scala 19:72:@10825.4]
  assign _T_26660 = _T_26659 | _T_26637; // @[Mux.scala 19:72:@10826.4]
  assign _T_26661 = _T_26660 | _T_26646; // @[Mux.scala 19:72:@10827.4]
  assign _T_26662 = _T_26661 | _T_26655; // @[Mux.scala 19:72:@10828.4]
  assign outputPriorityPorts_0_0 = _T_26662[0]; // @[Mux.scala 19:72:@10832.4]
  assign outputPriorityPorts_0_1 = _T_26662[1]; // @[Mux.scala 19:72:@10834.4]
  assign outputPriorityPorts_0_2 = _T_26662[2]; // @[Mux.scala 19:72:@10836.4]
  assign outputPriorityPorts_0_3 = _T_26662[3]; // @[Mux.scala 19:72:@10838.4]
  assign outputPriorityPorts_0_4 = _T_26662[4]; // @[Mux.scala 19:72:@10840.4]
  assign outputPriorityPorts_0_5 = _T_26662[5]; // @[Mux.scala 19:72:@10842.4]
  assign outputPriorityPorts_0_6 = _T_26662[6]; // @[Mux.scala 19:72:@10844.4]
  assign outputPriorityPorts_0_7 = _T_26662[7]; // @[Mux.scala 19:72:@10846.4]
  assign _T_26742 = portQ_0 & _T_25659; // @[LoadQueue.scala 298:83:@10857.4]
  assign _T_26745 = portQ_1 & _T_25662; // @[LoadQueue.scala 298:83:@10859.4]
  assign _T_26748 = portQ_2 & _T_25665; // @[LoadQueue.scala 298:83:@10861.4]
  assign _T_26751 = portQ_3 & _T_25668; // @[LoadQueue.scala 298:83:@10863.4]
  assign _T_26754 = portQ_4 & _T_25671; // @[LoadQueue.scala 298:83:@10865.4]
  assign _T_26757 = portQ_5 & _T_25674; // @[LoadQueue.scala 298:83:@10867.4]
  assign _T_26760 = portQ_6 & _T_25677; // @[LoadQueue.scala 298:83:@10869.4]
  assign _T_26763 = portQ_7 & _T_25680; // @[LoadQueue.scala 298:83:@10871.4]
  assign _T_26814 = _T_26763 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10901.4]
  assign _T_26815 = _T_26760 ? 8'h40 : _T_26814; // @[Mux.scala 31:69:@10902.4]
  assign _T_26816 = _T_26757 ? 8'h20 : _T_26815; // @[Mux.scala 31:69:@10903.4]
  assign _T_26817 = _T_26754 ? 8'h10 : _T_26816; // @[Mux.scala 31:69:@10904.4]
  assign _T_26818 = _T_26751 ? 8'h8 : _T_26817; // @[Mux.scala 31:69:@10905.4]
  assign _T_26819 = _T_26748 ? 8'h4 : _T_26818; // @[Mux.scala 31:69:@10906.4]
  assign _T_26820 = _T_26745 ? 8'h2 : _T_26819; // @[Mux.scala 31:69:@10907.4]
  assign _T_26821 = _T_26742 ? 8'h1 : _T_26820; // @[Mux.scala 31:69:@10908.4]
  assign _T_26822 = _T_26821[0]; // @[OneHot.scala 66:30:@10909.4]
  assign _T_26823 = _T_26821[1]; // @[OneHot.scala 66:30:@10910.4]
  assign _T_26824 = _T_26821[2]; // @[OneHot.scala 66:30:@10911.4]
  assign _T_26825 = _T_26821[3]; // @[OneHot.scala 66:30:@10912.4]
  assign _T_26826 = _T_26821[4]; // @[OneHot.scala 66:30:@10913.4]
  assign _T_26827 = _T_26821[5]; // @[OneHot.scala 66:30:@10914.4]
  assign _T_26828 = _T_26821[6]; // @[OneHot.scala 66:30:@10915.4]
  assign _T_26829 = _T_26821[7]; // @[OneHot.scala 66:30:@10916.4]
  assign _T_26854 = _T_26742 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10926.4]
  assign _T_26855 = _T_26763 ? 8'h40 : _T_26854; // @[Mux.scala 31:69:@10927.4]
  assign _T_26856 = _T_26760 ? 8'h20 : _T_26855; // @[Mux.scala 31:69:@10928.4]
  assign _T_26857 = _T_26757 ? 8'h10 : _T_26856; // @[Mux.scala 31:69:@10929.4]
  assign _T_26858 = _T_26754 ? 8'h8 : _T_26857; // @[Mux.scala 31:69:@10930.4]
  assign _T_26859 = _T_26751 ? 8'h4 : _T_26858; // @[Mux.scala 31:69:@10931.4]
  assign _T_26860 = _T_26748 ? 8'h2 : _T_26859; // @[Mux.scala 31:69:@10932.4]
  assign _T_26861 = _T_26745 ? 8'h1 : _T_26860; // @[Mux.scala 31:69:@10933.4]
  assign _T_26862 = _T_26861[0]; // @[OneHot.scala 66:30:@10934.4]
  assign _T_26863 = _T_26861[1]; // @[OneHot.scala 66:30:@10935.4]
  assign _T_26864 = _T_26861[2]; // @[OneHot.scala 66:30:@10936.4]
  assign _T_26865 = _T_26861[3]; // @[OneHot.scala 66:30:@10937.4]
  assign _T_26866 = _T_26861[4]; // @[OneHot.scala 66:30:@10938.4]
  assign _T_26867 = _T_26861[5]; // @[OneHot.scala 66:30:@10939.4]
  assign _T_26868 = _T_26861[6]; // @[OneHot.scala 66:30:@10940.4]
  assign _T_26869 = _T_26861[7]; // @[OneHot.scala 66:30:@10941.4]
  assign _T_26894 = _T_26745 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10951.4]
  assign _T_26895 = _T_26742 ? 8'h40 : _T_26894; // @[Mux.scala 31:69:@10952.4]
  assign _T_26896 = _T_26763 ? 8'h20 : _T_26895; // @[Mux.scala 31:69:@10953.4]
  assign _T_26897 = _T_26760 ? 8'h10 : _T_26896; // @[Mux.scala 31:69:@10954.4]
  assign _T_26898 = _T_26757 ? 8'h8 : _T_26897; // @[Mux.scala 31:69:@10955.4]
  assign _T_26899 = _T_26754 ? 8'h4 : _T_26898; // @[Mux.scala 31:69:@10956.4]
  assign _T_26900 = _T_26751 ? 8'h2 : _T_26899; // @[Mux.scala 31:69:@10957.4]
  assign _T_26901 = _T_26748 ? 8'h1 : _T_26900; // @[Mux.scala 31:69:@10958.4]
  assign _T_26902 = _T_26901[0]; // @[OneHot.scala 66:30:@10959.4]
  assign _T_26903 = _T_26901[1]; // @[OneHot.scala 66:30:@10960.4]
  assign _T_26904 = _T_26901[2]; // @[OneHot.scala 66:30:@10961.4]
  assign _T_26905 = _T_26901[3]; // @[OneHot.scala 66:30:@10962.4]
  assign _T_26906 = _T_26901[4]; // @[OneHot.scala 66:30:@10963.4]
  assign _T_26907 = _T_26901[5]; // @[OneHot.scala 66:30:@10964.4]
  assign _T_26908 = _T_26901[6]; // @[OneHot.scala 66:30:@10965.4]
  assign _T_26909 = _T_26901[7]; // @[OneHot.scala 66:30:@10966.4]
  assign _T_26934 = _T_26748 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@10976.4]
  assign _T_26935 = _T_26745 ? 8'h40 : _T_26934; // @[Mux.scala 31:69:@10977.4]
  assign _T_26936 = _T_26742 ? 8'h20 : _T_26935; // @[Mux.scala 31:69:@10978.4]
  assign _T_26937 = _T_26763 ? 8'h10 : _T_26936; // @[Mux.scala 31:69:@10979.4]
  assign _T_26938 = _T_26760 ? 8'h8 : _T_26937; // @[Mux.scala 31:69:@10980.4]
  assign _T_26939 = _T_26757 ? 8'h4 : _T_26938; // @[Mux.scala 31:69:@10981.4]
  assign _T_26940 = _T_26754 ? 8'h2 : _T_26939; // @[Mux.scala 31:69:@10982.4]
  assign _T_26941 = _T_26751 ? 8'h1 : _T_26940; // @[Mux.scala 31:69:@10983.4]
  assign _T_26942 = _T_26941[0]; // @[OneHot.scala 66:30:@10984.4]
  assign _T_26943 = _T_26941[1]; // @[OneHot.scala 66:30:@10985.4]
  assign _T_26944 = _T_26941[2]; // @[OneHot.scala 66:30:@10986.4]
  assign _T_26945 = _T_26941[3]; // @[OneHot.scala 66:30:@10987.4]
  assign _T_26946 = _T_26941[4]; // @[OneHot.scala 66:30:@10988.4]
  assign _T_26947 = _T_26941[5]; // @[OneHot.scala 66:30:@10989.4]
  assign _T_26948 = _T_26941[6]; // @[OneHot.scala 66:30:@10990.4]
  assign _T_26949 = _T_26941[7]; // @[OneHot.scala 66:30:@10991.4]
  assign _T_26974 = _T_26751 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11001.4]
  assign _T_26975 = _T_26748 ? 8'h40 : _T_26974; // @[Mux.scala 31:69:@11002.4]
  assign _T_26976 = _T_26745 ? 8'h20 : _T_26975; // @[Mux.scala 31:69:@11003.4]
  assign _T_26977 = _T_26742 ? 8'h10 : _T_26976; // @[Mux.scala 31:69:@11004.4]
  assign _T_26978 = _T_26763 ? 8'h8 : _T_26977; // @[Mux.scala 31:69:@11005.4]
  assign _T_26979 = _T_26760 ? 8'h4 : _T_26978; // @[Mux.scala 31:69:@11006.4]
  assign _T_26980 = _T_26757 ? 8'h2 : _T_26979; // @[Mux.scala 31:69:@11007.4]
  assign _T_26981 = _T_26754 ? 8'h1 : _T_26980; // @[Mux.scala 31:69:@11008.4]
  assign _T_26982 = _T_26981[0]; // @[OneHot.scala 66:30:@11009.4]
  assign _T_26983 = _T_26981[1]; // @[OneHot.scala 66:30:@11010.4]
  assign _T_26984 = _T_26981[2]; // @[OneHot.scala 66:30:@11011.4]
  assign _T_26985 = _T_26981[3]; // @[OneHot.scala 66:30:@11012.4]
  assign _T_26986 = _T_26981[4]; // @[OneHot.scala 66:30:@11013.4]
  assign _T_26987 = _T_26981[5]; // @[OneHot.scala 66:30:@11014.4]
  assign _T_26988 = _T_26981[6]; // @[OneHot.scala 66:30:@11015.4]
  assign _T_26989 = _T_26981[7]; // @[OneHot.scala 66:30:@11016.4]
  assign _T_27014 = _T_26754 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11026.4]
  assign _T_27015 = _T_26751 ? 8'h40 : _T_27014; // @[Mux.scala 31:69:@11027.4]
  assign _T_27016 = _T_26748 ? 8'h20 : _T_27015; // @[Mux.scala 31:69:@11028.4]
  assign _T_27017 = _T_26745 ? 8'h10 : _T_27016; // @[Mux.scala 31:69:@11029.4]
  assign _T_27018 = _T_26742 ? 8'h8 : _T_27017; // @[Mux.scala 31:69:@11030.4]
  assign _T_27019 = _T_26763 ? 8'h4 : _T_27018; // @[Mux.scala 31:69:@11031.4]
  assign _T_27020 = _T_26760 ? 8'h2 : _T_27019; // @[Mux.scala 31:69:@11032.4]
  assign _T_27021 = _T_26757 ? 8'h1 : _T_27020; // @[Mux.scala 31:69:@11033.4]
  assign _T_27022 = _T_27021[0]; // @[OneHot.scala 66:30:@11034.4]
  assign _T_27023 = _T_27021[1]; // @[OneHot.scala 66:30:@11035.4]
  assign _T_27024 = _T_27021[2]; // @[OneHot.scala 66:30:@11036.4]
  assign _T_27025 = _T_27021[3]; // @[OneHot.scala 66:30:@11037.4]
  assign _T_27026 = _T_27021[4]; // @[OneHot.scala 66:30:@11038.4]
  assign _T_27027 = _T_27021[5]; // @[OneHot.scala 66:30:@11039.4]
  assign _T_27028 = _T_27021[6]; // @[OneHot.scala 66:30:@11040.4]
  assign _T_27029 = _T_27021[7]; // @[OneHot.scala 66:30:@11041.4]
  assign _T_27054 = _T_26757 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11051.4]
  assign _T_27055 = _T_26754 ? 8'h40 : _T_27054; // @[Mux.scala 31:69:@11052.4]
  assign _T_27056 = _T_26751 ? 8'h20 : _T_27055; // @[Mux.scala 31:69:@11053.4]
  assign _T_27057 = _T_26748 ? 8'h10 : _T_27056; // @[Mux.scala 31:69:@11054.4]
  assign _T_27058 = _T_26745 ? 8'h8 : _T_27057; // @[Mux.scala 31:69:@11055.4]
  assign _T_27059 = _T_26742 ? 8'h4 : _T_27058; // @[Mux.scala 31:69:@11056.4]
  assign _T_27060 = _T_26763 ? 8'h2 : _T_27059; // @[Mux.scala 31:69:@11057.4]
  assign _T_27061 = _T_26760 ? 8'h1 : _T_27060; // @[Mux.scala 31:69:@11058.4]
  assign _T_27062 = _T_27061[0]; // @[OneHot.scala 66:30:@11059.4]
  assign _T_27063 = _T_27061[1]; // @[OneHot.scala 66:30:@11060.4]
  assign _T_27064 = _T_27061[2]; // @[OneHot.scala 66:30:@11061.4]
  assign _T_27065 = _T_27061[3]; // @[OneHot.scala 66:30:@11062.4]
  assign _T_27066 = _T_27061[4]; // @[OneHot.scala 66:30:@11063.4]
  assign _T_27067 = _T_27061[5]; // @[OneHot.scala 66:30:@11064.4]
  assign _T_27068 = _T_27061[6]; // @[OneHot.scala 66:30:@11065.4]
  assign _T_27069 = _T_27061[7]; // @[OneHot.scala 66:30:@11066.4]
  assign _T_27094 = _T_26760 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11076.4]
  assign _T_27095 = _T_26757 ? 8'h40 : _T_27094; // @[Mux.scala 31:69:@11077.4]
  assign _T_27096 = _T_26754 ? 8'h20 : _T_27095; // @[Mux.scala 31:69:@11078.4]
  assign _T_27097 = _T_26751 ? 8'h10 : _T_27096; // @[Mux.scala 31:69:@11079.4]
  assign _T_27098 = _T_26748 ? 8'h8 : _T_27097; // @[Mux.scala 31:69:@11080.4]
  assign _T_27099 = _T_26745 ? 8'h4 : _T_27098; // @[Mux.scala 31:69:@11081.4]
  assign _T_27100 = _T_26742 ? 8'h2 : _T_27099; // @[Mux.scala 31:69:@11082.4]
  assign _T_27101 = _T_26763 ? 8'h1 : _T_27100; // @[Mux.scala 31:69:@11083.4]
  assign _T_27102 = _T_27101[0]; // @[OneHot.scala 66:30:@11084.4]
  assign _T_27103 = _T_27101[1]; // @[OneHot.scala 66:30:@11085.4]
  assign _T_27104 = _T_27101[2]; // @[OneHot.scala 66:30:@11086.4]
  assign _T_27105 = _T_27101[3]; // @[OneHot.scala 66:30:@11087.4]
  assign _T_27106 = _T_27101[4]; // @[OneHot.scala 66:30:@11088.4]
  assign _T_27107 = _T_27101[5]; // @[OneHot.scala 66:30:@11089.4]
  assign _T_27108 = _T_27101[6]; // @[OneHot.scala 66:30:@11090.4]
  assign _T_27109 = _T_27101[7]; // @[OneHot.scala 66:30:@11091.4]
  assign _T_27150 = {_T_26829,_T_26828,_T_26827,_T_26826,_T_26825,_T_26824,_T_26823,_T_26822}; // @[Mux.scala 19:72:@11107.4]
  assign _T_27152 = _T_24152 ? _T_27150 : 8'h0; // @[Mux.scala 19:72:@11108.4]
  assign _T_27159 = {_T_26868,_T_26867,_T_26866,_T_26865,_T_26864,_T_26863,_T_26862,_T_26869}; // @[Mux.scala 19:72:@11115.4]
  assign _T_27161 = _T_24153 ? _T_27159 : 8'h0; // @[Mux.scala 19:72:@11116.4]
  assign _T_27168 = {_T_26907,_T_26906,_T_26905,_T_26904,_T_26903,_T_26902,_T_26909,_T_26908}; // @[Mux.scala 19:72:@11123.4]
  assign _T_27170 = _T_24154 ? _T_27168 : 8'h0; // @[Mux.scala 19:72:@11124.4]
  assign _T_27177 = {_T_26946,_T_26945,_T_26944,_T_26943,_T_26942,_T_26949,_T_26948,_T_26947}; // @[Mux.scala 19:72:@11131.4]
  assign _T_27179 = _T_24155 ? _T_27177 : 8'h0; // @[Mux.scala 19:72:@11132.4]
  assign _T_27186 = {_T_26985,_T_26984,_T_26983,_T_26982,_T_26989,_T_26988,_T_26987,_T_26986}; // @[Mux.scala 19:72:@11139.4]
  assign _T_27188 = _T_24156 ? _T_27186 : 8'h0; // @[Mux.scala 19:72:@11140.4]
  assign _T_27195 = {_T_27024,_T_27023,_T_27022,_T_27029,_T_27028,_T_27027,_T_27026,_T_27025}; // @[Mux.scala 19:72:@11147.4]
  assign _T_27197 = _T_24157 ? _T_27195 : 8'h0; // @[Mux.scala 19:72:@11148.4]
  assign _T_27204 = {_T_27063,_T_27062,_T_27069,_T_27068,_T_27067,_T_27066,_T_27065,_T_27064}; // @[Mux.scala 19:72:@11155.4]
  assign _T_27206 = _T_24158 ? _T_27204 : 8'h0; // @[Mux.scala 19:72:@11156.4]
  assign _T_27213 = {_T_27102,_T_27109,_T_27108,_T_27107,_T_27106,_T_27105,_T_27104,_T_27103}; // @[Mux.scala 19:72:@11163.4]
  assign _T_27215 = _T_24159 ? _T_27213 : 8'h0; // @[Mux.scala 19:72:@11164.4]
  assign _T_27216 = _T_27152 | _T_27161; // @[Mux.scala 19:72:@11165.4]
  assign _T_27217 = _T_27216 | _T_27170; // @[Mux.scala 19:72:@11166.4]
  assign _T_27218 = _T_27217 | _T_27179; // @[Mux.scala 19:72:@11167.4]
  assign _T_27219 = _T_27218 | _T_27188; // @[Mux.scala 19:72:@11168.4]
  assign _T_27220 = _T_27219 | _T_27197; // @[Mux.scala 19:72:@11169.4]
  assign _T_27221 = _T_27220 | _T_27206; // @[Mux.scala 19:72:@11170.4]
  assign _T_27222 = _T_27221 | _T_27215; // @[Mux.scala 19:72:@11171.4]
  assign inputPriorityPorts_1_0 = _T_27222[0]; // @[Mux.scala 19:72:@11175.4]
  assign inputPriorityPorts_1_1 = _T_27222[1]; // @[Mux.scala 19:72:@11177.4]
  assign inputPriorityPorts_1_2 = _T_27222[2]; // @[Mux.scala 19:72:@11179.4]
  assign inputPriorityPorts_1_3 = _T_27222[3]; // @[Mux.scala 19:72:@11181.4]
  assign inputPriorityPorts_1_4 = _T_27222[4]; // @[Mux.scala 19:72:@11183.4]
  assign inputPriorityPorts_1_5 = _T_27222[5]; // @[Mux.scala 19:72:@11185.4]
  assign inputPriorityPorts_1_6 = _T_27222[6]; // @[Mux.scala 19:72:@11187.4]
  assign inputPriorityPorts_1_7 = _T_27222[7]; // @[Mux.scala 19:72:@11189.4]
  assign _T_27336 = portQ_7 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11219.4]
  assign _T_27337 = portQ_6 ? 8'h40 : _T_27336; // @[Mux.scala 31:69:@11220.4]
  assign _T_27338 = portQ_5 ? 8'h20 : _T_27337; // @[Mux.scala 31:69:@11221.4]
  assign _T_27339 = portQ_4 ? 8'h10 : _T_27338; // @[Mux.scala 31:69:@11222.4]
  assign _T_27340 = portQ_3 ? 8'h8 : _T_27339; // @[Mux.scala 31:69:@11223.4]
  assign _T_27341 = portQ_2 ? 8'h4 : _T_27340; // @[Mux.scala 31:69:@11224.4]
  assign _T_27342 = portQ_1 ? 8'h2 : _T_27341; // @[Mux.scala 31:69:@11225.4]
  assign _T_27343 = portQ_0 ? 8'h1 : _T_27342; // @[Mux.scala 31:69:@11226.4]
  assign _T_27344 = _T_27343[0]; // @[OneHot.scala 66:30:@11227.4]
  assign _T_27345 = _T_27343[1]; // @[OneHot.scala 66:30:@11228.4]
  assign _T_27346 = _T_27343[2]; // @[OneHot.scala 66:30:@11229.4]
  assign _T_27347 = _T_27343[3]; // @[OneHot.scala 66:30:@11230.4]
  assign _T_27348 = _T_27343[4]; // @[OneHot.scala 66:30:@11231.4]
  assign _T_27349 = _T_27343[5]; // @[OneHot.scala 66:30:@11232.4]
  assign _T_27350 = _T_27343[6]; // @[OneHot.scala 66:30:@11233.4]
  assign _T_27351 = _T_27343[7]; // @[OneHot.scala 66:30:@11234.4]
  assign _T_27376 = portQ_0 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11244.4]
  assign _T_27377 = portQ_7 ? 8'h40 : _T_27376; // @[Mux.scala 31:69:@11245.4]
  assign _T_27378 = portQ_6 ? 8'h20 : _T_27377; // @[Mux.scala 31:69:@11246.4]
  assign _T_27379 = portQ_5 ? 8'h10 : _T_27378; // @[Mux.scala 31:69:@11247.4]
  assign _T_27380 = portQ_4 ? 8'h8 : _T_27379; // @[Mux.scala 31:69:@11248.4]
  assign _T_27381 = portQ_3 ? 8'h4 : _T_27380; // @[Mux.scala 31:69:@11249.4]
  assign _T_27382 = portQ_2 ? 8'h2 : _T_27381; // @[Mux.scala 31:69:@11250.4]
  assign _T_27383 = portQ_1 ? 8'h1 : _T_27382; // @[Mux.scala 31:69:@11251.4]
  assign _T_27384 = _T_27383[0]; // @[OneHot.scala 66:30:@11252.4]
  assign _T_27385 = _T_27383[1]; // @[OneHot.scala 66:30:@11253.4]
  assign _T_27386 = _T_27383[2]; // @[OneHot.scala 66:30:@11254.4]
  assign _T_27387 = _T_27383[3]; // @[OneHot.scala 66:30:@11255.4]
  assign _T_27388 = _T_27383[4]; // @[OneHot.scala 66:30:@11256.4]
  assign _T_27389 = _T_27383[5]; // @[OneHot.scala 66:30:@11257.4]
  assign _T_27390 = _T_27383[6]; // @[OneHot.scala 66:30:@11258.4]
  assign _T_27391 = _T_27383[7]; // @[OneHot.scala 66:30:@11259.4]
  assign _T_27416 = portQ_1 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11269.4]
  assign _T_27417 = portQ_0 ? 8'h40 : _T_27416; // @[Mux.scala 31:69:@11270.4]
  assign _T_27418 = portQ_7 ? 8'h20 : _T_27417; // @[Mux.scala 31:69:@11271.4]
  assign _T_27419 = portQ_6 ? 8'h10 : _T_27418; // @[Mux.scala 31:69:@11272.4]
  assign _T_27420 = portQ_5 ? 8'h8 : _T_27419; // @[Mux.scala 31:69:@11273.4]
  assign _T_27421 = portQ_4 ? 8'h4 : _T_27420; // @[Mux.scala 31:69:@11274.4]
  assign _T_27422 = portQ_3 ? 8'h2 : _T_27421; // @[Mux.scala 31:69:@11275.4]
  assign _T_27423 = portQ_2 ? 8'h1 : _T_27422; // @[Mux.scala 31:69:@11276.4]
  assign _T_27424 = _T_27423[0]; // @[OneHot.scala 66:30:@11277.4]
  assign _T_27425 = _T_27423[1]; // @[OneHot.scala 66:30:@11278.4]
  assign _T_27426 = _T_27423[2]; // @[OneHot.scala 66:30:@11279.4]
  assign _T_27427 = _T_27423[3]; // @[OneHot.scala 66:30:@11280.4]
  assign _T_27428 = _T_27423[4]; // @[OneHot.scala 66:30:@11281.4]
  assign _T_27429 = _T_27423[5]; // @[OneHot.scala 66:30:@11282.4]
  assign _T_27430 = _T_27423[6]; // @[OneHot.scala 66:30:@11283.4]
  assign _T_27431 = _T_27423[7]; // @[OneHot.scala 66:30:@11284.4]
  assign _T_27456 = portQ_2 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11294.4]
  assign _T_27457 = portQ_1 ? 8'h40 : _T_27456; // @[Mux.scala 31:69:@11295.4]
  assign _T_27458 = portQ_0 ? 8'h20 : _T_27457; // @[Mux.scala 31:69:@11296.4]
  assign _T_27459 = portQ_7 ? 8'h10 : _T_27458; // @[Mux.scala 31:69:@11297.4]
  assign _T_27460 = portQ_6 ? 8'h8 : _T_27459; // @[Mux.scala 31:69:@11298.4]
  assign _T_27461 = portQ_5 ? 8'h4 : _T_27460; // @[Mux.scala 31:69:@11299.4]
  assign _T_27462 = portQ_4 ? 8'h2 : _T_27461; // @[Mux.scala 31:69:@11300.4]
  assign _T_27463 = portQ_3 ? 8'h1 : _T_27462; // @[Mux.scala 31:69:@11301.4]
  assign _T_27464 = _T_27463[0]; // @[OneHot.scala 66:30:@11302.4]
  assign _T_27465 = _T_27463[1]; // @[OneHot.scala 66:30:@11303.4]
  assign _T_27466 = _T_27463[2]; // @[OneHot.scala 66:30:@11304.4]
  assign _T_27467 = _T_27463[3]; // @[OneHot.scala 66:30:@11305.4]
  assign _T_27468 = _T_27463[4]; // @[OneHot.scala 66:30:@11306.4]
  assign _T_27469 = _T_27463[5]; // @[OneHot.scala 66:30:@11307.4]
  assign _T_27470 = _T_27463[6]; // @[OneHot.scala 66:30:@11308.4]
  assign _T_27471 = _T_27463[7]; // @[OneHot.scala 66:30:@11309.4]
  assign _T_27496 = portQ_3 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11319.4]
  assign _T_27497 = portQ_2 ? 8'h40 : _T_27496; // @[Mux.scala 31:69:@11320.4]
  assign _T_27498 = portQ_1 ? 8'h20 : _T_27497; // @[Mux.scala 31:69:@11321.4]
  assign _T_27499 = portQ_0 ? 8'h10 : _T_27498; // @[Mux.scala 31:69:@11322.4]
  assign _T_27500 = portQ_7 ? 8'h8 : _T_27499; // @[Mux.scala 31:69:@11323.4]
  assign _T_27501 = portQ_6 ? 8'h4 : _T_27500; // @[Mux.scala 31:69:@11324.4]
  assign _T_27502 = portQ_5 ? 8'h2 : _T_27501; // @[Mux.scala 31:69:@11325.4]
  assign _T_27503 = portQ_4 ? 8'h1 : _T_27502; // @[Mux.scala 31:69:@11326.4]
  assign _T_27504 = _T_27503[0]; // @[OneHot.scala 66:30:@11327.4]
  assign _T_27505 = _T_27503[1]; // @[OneHot.scala 66:30:@11328.4]
  assign _T_27506 = _T_27503[2]; // @[OneHot.scala 66:30:@11329.4]
  assign _T_27507 = _T_27503[3]; // @[OneHot.scala 66:30:@11330.4]
  assign _T_27508 = _T_27503[4]; // @[OneHot.scala 66:30:@11331.4]
  assign _T_27509 = _T_27503[5]; // @[OneHot.scala 66:30:@11332.4]
  assign _T_27510 = _T_27503[6]; // @[OneHot.scala 66:30:@11333.4]
  assign _T_27511 = _T_27503[7]; // @[OneHot.scala 66:30:@11334.4]
  assign _T_27536 = portQ_4 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11344.4]
  assign _T_27537 = portQ_3 ? 8'h40 : _T_27536; // @[Mux.scala 31:69:@11345.4]
  assign _T_27538 = portQ_2 ? 8'h20 : _T_27537; // @[Mux.scala 31:69:@11346.4]
  assign _T_27539 = portQ_1 ? 8'h10 : _T_27538; // @[Mux.scala 31:69:@11347.4]
  assign _T_27540 = portQ_0 ? 8'h8 : _T_27539; // @[Mux.scala 31:69:@11348.4]
  assign _T_27541 = portQ_7 ? 8'h4 : _T_27540; // @[Mux.scala 31:69:@11349.4]
  assign _T_27542 = portQ_6 ? 8'h2 : _T_27541; // @[Mux.scala 31:69:@11350.4]
  assign _T_27543 = portQ_5 ? 8'h1 : _T_27542; // @[Mux.scala 31:69:@11351.4]
  assign _T_27544 = _T_27543[0]; // @[OneHot.scala 66:30:@11352.4]
  assign _T_27545 = _T_27543[1]; // @[OneHot.scala 66:30:@11353.4]
  assign _T_27546 = _T_27543[2]; // @[OneHot.scala 66:30:@11354.4]
  assign _T_27547 = _T_27543[3]; // @[OneHot.scala 66:30:@11355.4]
  assign _T_27548 = _T_27543[4]; // @[OneHot.scala 66:30:@11356.4]
  assign _T_27549 = _T_27543[5]; // @[OneHot.scala 66:30:@11357.4]
  assign _T_27550 = _T_27543[6]; // @[OneHot.scala 66:30:@11358.4]
  assign _T_27551 = _T_27543[7]; // @[OneHot.scala 66:30:@11359.4]
  assign _T_27576 = portQ_5 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11369.4]
  assign _T_27577 = portQ_4 ? 8'h40 : _T_27576; // @[Mux.scala 31:69:@11370.4]
  assign _T_27578 = portQ_3 ? 8'h20 : _T_27577; // @[Mux.scala 31:69:@11371.4]
  assign _T_27579 = portQ_2 ? 8'h10 : _T_27578; // @[Mux.scala 31:69:@11372.4]
  assign _T_27580 = portQ_1 ? 8'h8 : _T_27579; // @[Mux.scala 31:69:@11373.4]
  assign _T_27581 = portQ_0 ? 8'h4 : _T_27580; // @[Mux.scala 31:69:@11374.4]
  assign _T_27582 = portQ_7 ? 8'h2 : _T_27581; // @[Mux.scala 31:69:@11375.4]
  assign _T_27583 = portQ_6 ? 8'h1 : _T_27582; // @[Mux.scala 31:69:@11376.4]
  assign _T_27584 = _T_27583[0]; // @[OneHot.scala 66:30:@11377.4]
  assign _T_27585 = _T_27583[1]; // @[OneHot.scala 66:30:@11378.4]
  assign _T_27586 = _T_27583[2]; // @[OneHot.scala 66:30:@11379.4]
  assign _T_27587 = _T_27583[3]; // @[OneHot.scala 66:30:@11380.4]
  assign _T_27588 = _T_27583[4]; // @[OneHot.scala 66:30:@11381.4]
  assign _T_27589 = _T_27583[5]; // @[OneHot.scala 66:30:@11382.4]
  assign _T_27590 = _T_27583[6]; // @[OneHot.scala 66:30:@11383.4]
  assign _T_27591 = _T_27583[7]; // @[OneHot.scala 66:30:@11384.4]
  assign _T_27616 = portQ_6 ? 8'h80 : 8'h0; // @[Mux.scala 31:69:@11394.4]
  assign _T_27617 = portQ_5 ? 8'h40 : _T_27616; // @[Mux.scala 31:69:@11395.4]
  assign _T_27618 = portQ_4 ? 8'h20 : _T_27617; // @[Mux.scala 31:69:@11396.4]
  assign _T_27619 = portQ_3 ? 8'h10 : _T_27618; // @[Mux.scala 31:69:@11397.4]
  assign _T_27620 = portQ_2 ? 8'h8 : _T_27619; // @[Mux.scala 31:69:@11398.4]
  assign _T_27621 = portQ_1 ? 8'h4 : _T_27620; // @[Mux.scala 31:69:@11399.4]
  assign _T_27622 = portQ_0 ? 8'h2 : _T_27621; // @[Mux.scala 31:69:@11400.4]
  assign _T_27623 = portQ_7 ? 8'h1 : _T_27622; // @[Mux.scala 31:69:@11401.4]
  assign _T_27624 = _T_27623[0]; // @[OneHot.scala 66:30:@11402.4]
  assign _T_27625 = _T_27623[1]; // @[OneHot.scala 66:30:@11403.4]
  assign _T_27626 = _T_27623[2]; // @[OneHot.scala 66:30:@11404.4]
  assign _T_27627 = _T_27623[3]; // @[OneHot.scala 66:30:@11405.4]
  assign _T_27628 = _T_27623[4]; // @[OneHot.scala 66:30:@11406.4]
  assign _T_27629 = _T_27623[5]; // @[OneHot.scala 66:30:@11407.4]
  assign _T_27630 = _T_27623[6]; // @[OneHot.scala 66:30:@11408.4]
  assign _T_27631 = _T_27623[7]; // @[OneHot.scala 66:30:@11409.4]
  assign _T_27672 = {_T_27351,_T_27350,_T_27349,_T_27348,_T_27347,_T_27346,_T_27345,_T_27344}; // @[Mux.scala 19:72:@11425.4]
  assign _T_27674 = _T_24152 ? _T_27672 : 8'h0; // @[Mux.scala 19:72:@11426.4]
  assign _T_27681 = {_T_27390,_T_27389,_T_27388,_T_27387,_T_27386,_T_27385,_T_27384,_T_27391}; // @[Mux.scala 19:72:@11433.4]
  assign _T_27683 = _T_24153 ? _T_27681 : 8'h0; // @[Mux.scala 19:72:@11434.4]
  assign _T_27690 = {_T_27429,_T_27428,_T_27427,_T_27426,_T_27425,_T_27424,_T_27431,_T_27430}; // @[Mux.scala 19:72:@11441.4]
  assign _T_27692 = _T_24154 ? _T_27690 : 8'h0; // @[Mux.scala 19:72:@11442.4]
  assign _T_27699 = {_T_27468,_T_27467,_T_27466,_T_27465,_T_27464,_T_27471,_T_27470,_T_27469}; // @[Mux.scala 19:72:@11449.4]
  assign _T_27701 = _T_24155 ? _T_27699 : 8'h0; // @[Mux.scala 19:72:@11450.4]
  assign _T_27708 = {_T_27507,_T_27506,_T_27505,_T_27504,_T_27511,_T_27510,_T_27509,_T_27508}; // @[Mux.scala 19:72:@11457.4]
  assign _T_27710 = _T_24156 ? _T_27708 : 8'h0; // @[Mux.scala 19:72:@11458.4]
  assign _T_27717 = {_T_27546,_T_27545,_T_27544,_T_27551,_T_27550,_T_27549,_T_27548,_T_27547}; // @[Mux.scala 19:72:@11465.4]
  assign _T_27719 = _T_24157 ? _T_27717 : 8'h0; // @[Mux.scala 19:72:@11466.4]
  assign _T_27726 = {_T_27585,_T_27584,_T_27591,_T_27590,_T_27589,_T_27588,_T_27587,_T_27586}; // @[Mux.scala 19:72:@11473.4]
  assign _T_27728 = _T_24158 ? _T_27726 : 8'h0; // @[Mux.scala 19:72:@11474.4]
  assign _T_27735 = {_T_27624,_T_27631,_T_27630,_T_27629,_T_27628,_T_27627,_T_27626,_T_27625}; // @[Mux.scala 19:72:@11481.4]
  assign _T_27737 = _T_24159 ? _T_27735 : 8'h0; // @[Mux.scala 19:72:@11482.4]
  assign _T_27738 = _T_27674 | _T_27683; // @[Mux.scala 19:72:@11483.4]
  assign _T_27739 = _T_27738 | _T_27692; // @[Mux.scala 19:72:@11484.4]
  assign _T_27740 = _T_27739 | _T_27701; // @[Mux.scala 19:72:@11485.4]
  assign _T_27741 = _T_27740 | _T_27710; // @[Mux.scala 19:72:@11486.4]
  assign _T_27742 = _T_27741 | _T_27719; // @[Mux.scala 19:72:@11487.4]
  assign _T_27743 = _T_27742 | _T_27728; // @[Mux.scala 19:72:@11488.4]
  assign _T_27744 = _T_27743 | _T_27737; // @[Mux.scala 19:72:@11489.4]
  assign outputPriorityPorts_1_0 = _T_27744[0]; // @[Mux.scala 19:72:@11493.4]
  assign outputPriorityPorts_1_1 = _T_27744[1]; // @[Mux.scala 19:72:@11495.4]
  assign outputPriorityPorts_1_2 = _T_27744[2]; // @[Mux.scala 19:72:@11497.4]
  assign outputPriorityPorts_1_3 = _T_27744[3]; // @[Mux.scala 19:72:@11499.4]
  assign outputPriorityPorts_1_4 = _T_27744[4]; // @[Mux.scala 19:72:@11501.4]
  assign outputPriorityPorts_1_5 = _T_27744[5]; // @[Mux.scala 19:72:@11503.4]
  assign outputPriorityPorts_1_6 = _T_27744[6]; // @[Mux.scala 19:72:@11505.4]
  assign outputPriorityPorts_1_7 = _T_27744[7]; // @[Mux.scala 19:72:@11507.4]
  assign _T_27823 = inputPriorityPorts_0_0 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@11521.6]
  assign _T_27824 = inputPriorityPorts_1_0 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@11522.6]
  assign _T_27835 = _T_27823 | _T_27824; // @[LoadQueue.scala 314:26:@11527.6]
  assign _T_27836 = {_T_27824,_T_27823}; // @[OneHot.scala 18:45:@11529.8]
  assign _T_27837 = _T_27836[1]; // @[CircuitMath.scala 30:8:@11530.8]
  assign _GEN_611 = _T_27837 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@11531.8]
  assign _GEN_612 = _T_27835 ? _GEN_611 : addrQ_0; // @[LoadQueue.scala 314:36:@11528.6]
  assign _GEN_613 = _T_27835 ? 1'h1 : addrKnown_0; // @[LoadQueue.scala 314:36:@11528.6]
  assign _GEN_614 = initBits_0 ? 1'h0 : _GEN_613; // @[LoadQueue.scala 308:34:@11517.4]
  assign _GEN_615 = initBits_0 ? addrQ_0 : _GEN_612; // @[LoadQueue.scala 308:34:@11517.4]
  assign _T_27841 = inputPriorityPorts_0_1 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@11539.6]
  assign _T_27842 = inputPriorityPorts_1_1 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@11540.6]
  assign _T_27853 = _T_27841 | _T_27842; // @[LoadQueue.scala 314:26:@11545.6]
  assign _T_27854 = {_T_27842,_T_27841}; // @[OneHot.scala 18:45:@11547.8]
  assign _T_27855 = _T_27854[1]; // @[CircuitMath.scala 30:8:@11548.8]
  assign _GEN_617 = _T_27855 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@11549.8]
  assign _GEN_618 = _T_27853 ? _GEN_617 : addrQ_1; // @[LoadQueue.scala 314:36:@11546.6]
  assign _GEN_619 = _T_27853 ? 1'h1 : addrKnown_1; // @[LoadQueue.scala 314:36:@11546.6]
  assign _GEN_620 = initBits_1 ? 1'h0 : _GEN_619; // @[LoadQueue.scala 308:34:@11535.4]
  assign _GEN_621 = initBits_1 ? addrQ_1 : _GEN_618; // @[LoadQueue.scala 308:34:@11535.4]
  assign _T_27859 = inputPriorityPorts_0_2 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@11557.6]
  assign _T_27860 = inputPriorityPorts_1_2 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@11558.6]
  assign _T_27871 = _T_27859 | _T_27860; // @[LoadQueue.scala 314:26:@11563.6]
  assign _T_27872 = {_T_27860,_T_27859}; // @[OneHot.scala 18:45:@11565.8]
  assign _T_27873 = _T_27872[1]; // @[CircuitMath.scala 30:8:@11566.8]
  assign _GEN_623 = _T_27873 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@11567.8]
  assign _GEN_624 = _T_27871 ? _GEN_623 : addrQ_2; // @[LoadQueue.scala 314:36:@11564.6]
  assign _GEN_625 = _T_27871 ? 1'h1 : addrKnown_2; // @[LoadQueue.scala 314:36:@11564.6]
  assign _GEN_626 = initBits_2 ? 1'h0 : _GEN_625; // @[LoadQueue.scala 308:34:@11553.4]
  assign _GEN_627 = initBits_2 ? addrQ_2 : _GEN_624; // @[LoadQueue.scala 308:34:@11553.4]
  assign _T_27877 = inputPriorityPorts_0_3 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@11575.6]
  assign _T_27878 = inputPriorityPorts_1_3 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@11576.6]
  assign _T_27889 = _T_27877 | _T_27878; // @[LoadQueue.scala 314:26:@11581.6]
  assign _T_27890 = {_T_27878,_T_27877}; // @[OneHot.scala 18:45:@11583.8]
  assign _T_27891 = _T_27890[1]; // @[CircuitMath.scala 30:8:@11584.8]
  assign _GEN_629 = _T_27891 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@11585.8]
  assign _GEN_630 = _T_27889 ? _GEN_629 : addrQ_3; // @[LoadQueue.scala 314:36:@11582.6]
  assign _GEN_631 = _T_27889 ? 1'h1 : addrKnown_3; // @[LoadQueue.scala 314:36:@11582.6]
  assign _GEN_632 = initBits_3 ? 1'h0 : _GEN_631; // @[LoadQueue.scala 308:34:@11571.4]
  assign _GEN_633 = initBits_3 ? addrQ_3 : _GEN_630; // @[LoadQueue.scala 308:34:@11571.4]
  assign _T_27895 = inputPriorityPorts_0_4 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@11593.6]
  assign _T_27896 = inputPriorityPorts_1_4 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@11594.6]
  assign _T_27907 = _T_27895 | _T_27896; // @[LoadQueue.scala 314:26:@11599.6]
  assign _T_27908 = {_T_27896,_T_27895}; // @[OneHot.scala 18:45:@11601.8]
  assign _T_27909 = _T_27908[1]; // @[CircuitMath.scala 30:8:@11602.8]
  assign _GEN_635 = _T_27909 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@11603.8]
  assign _GEN_636 = _T_27907 ? _GEN_635 : addrQ_4; // @[LoadQueue.scala 314:36:@11600.6]
  assign _GEN_637 = _T_27907 ? 1'h1 : addrKnown_4; // @[LoadQueue.scala 314:36:@11600.6]
  assign _GEN_638 = initBits_4 ? 1'h0 : _GEN_637; // @[LoadQueue.scala 308:34:@11589.4]
  assign _GEN_639 = initBits_4 ? addrQ_4 : _GEN_636; // @[LoadQueue.scala 308:34:@11589.4]
  assign _T_27913 = inputPriorityPorts_0_5 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@11611.6]
  assign _T_27914 = inputPriorityPorts_1_5 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@11612.6]
  assign _T_27925 = _T_27913 | _T_27914; // @[LoadQueue.scala 314:26:@11617.6]
  assign _T_27926 = {_T_27914,_T_27913}; // @[OneHot.scala 18:45:@11619.8]
  assign _T_27927 = _T_27926[1]; // @[CircuitMath.scala 30:8:@11620.8]
  assign _GEN_641 = _T_27927 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@11621.8]
  assign _GEN_642 = _T_27925 ? _GEN_641 : addrQ_5; // @[LoadQueue.scala 314:36:@11618.6]
  assign _GEN_643 = _T_27925 ? 1'h1 : addrKnown_5; // @[LoadQueue.scala 314:36:@11618.6]
  assign _GEN_644 = initBits_5 ? 1'h0 : _GEN_643; // @[LoadQueue.scala 308:34:@11607.4]
  assign _GEN_645 = initBits_5 ? addrQ_5 : _GEN_642; // @[LoadQueue.scala 308:34:@11607.4]
  assign _T_27931 = inputPriorityPorts_0_6 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@11629.6]
  assign _T_27932 = inputPriorityPorts_1_6 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@11630.6]
  assign _T_27943 = _T_27931 | _T_27932; // @[LoadQueue.scala 314:26:@11635.6]
  assign _T_27944 = {_T_27932,_T_27931}; // @[OneHot.scala 18:45:@11637.8]
  assign _T_27945 = _T_27944[1]; // @[CircuitMath.scala 30:8:@11638.8]
  assign _GEN_647 = _T_27945 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@11639.8]
  assign _GEN_648 = _T_27943 ? _GEN_647 : addrQ_6; // @[LoadQueue.scala 314:36:@11636.6]
  assign _GEN_649 = _T_27943 ? 1'h1 : addrKnown_6; // @[LoadQueue.scala 314:36:@11636.6]
  assign _GEN_650 = initBits_6 ? 1'h0 : _GEN_649; // @[LoadQueue.scala 308:34:@11625.4]
  assign _GEN_651 = initBits_6 ? addrQ_6 : _GEN_648; // @[LoadQueue.scala 308:34:@11625.4]
  assign _T_27949 = inputPriorityPorts_0_7 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@11647.6]
  assign _T_27950 = inputPriorityPorts_1_7 & io_loadAddrEnable_1; // @[LoadQueue.scala 313:47:@11648.6]
  assign _T_27961 = _T_27949 | _T_27950; // @[LoadQueue.scala 314:26:@11653.6]
  assign _T_27962 = {_T_27950,_T_27949}; // @[OneHot.scala 18:45:@11655.8]
  assign _T_27963 = _T_27962[1]; // @[CircuitMath.scala 30:8:@11656.8]
  assign _GEN_653 = _T_27963 ? io_addrFromLoadPorts_1 : io_addrFromLoadPorts_0; // @[LoadQueue.scala 315:29:@11657.8]
  assign _GEN_654 = _T_27961 ? _GEN_653 : addrQ_7; // @[LoadQueue.scala 314:36:@11654.6]
  assign _GEN_655 = _T_27961 ? 1'h1 : addrKnown_7; // @[LoadQueue.scala 314:36:@11654.6]
  assign _GEN_656 = initBits_7 ? 1'h0 : _GEN_655; // @[LoadQueue.scala 308:34:@11643.4]
  assign _GEN_657 = initBits_7 ? addrQ_7 : _GEN_654; // @[LoadQueue.scala 308:34:@11643.4]
  assign _T_27979 = outputPriorityPorts_0_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@11662.4]
  assign _T_27981 = loadCompleted_0 == 1'h0; // @[LoadQueue.scala 327:34:@11663.4]
  assign _T_27982 = _T_27979 & _T_27981; // @[LoadQueue.scala 327:31:@11664.4]
  assign _T_27983 = _T_27982 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@11665.4]
  assign _T_27984 = outputPriorityPorts_1_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@11666.4]
  assign _T_27987 = _T_27984 & _T_27981; // @[LoadQueue.scala 327:31:@11668.4]
  assign _T_27988 = _T_27987 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@11669.4]
  assign loadCompleting_0 = _T_27983 | _T_27988; // @[LoadQueue.scala 328:51:@11674.4]
  assign _T_28000 = outputPriorityPorts_0_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@11676.4]
  assign _T_28002 = loadCompleted_1 == 1'h0; // @[LoadQueue.scala 327:34:@11677.4]
  assign _T_28003 = _T_28000 & _T_28002; // @[LoadQueue.scala 327:31:@11678.4]
  assign _T_28004 = _T_28003 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@11679.4]
  assign _T_28005 = outputPriorityPorts_1_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@11680.4]
  assign _T_28008 = _T_28005 & _T_28002; // @[LoadQueue.scala 327:31:@11682.4]
  assign _T_28009 = _T_28008 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@11683.4]
  assign loadCompleting_1 = _T_28004 | _T_28009; // @[LoadQueue.scala 328:51:@11688.4]
  assign _T_28021 = outputPriorityPorts_0_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@11690.4]
  assign _T_28023 = loadCompleted_2 == 1'h0; // @[LoadQueue.scala 327:34:@11691.4]
  assign _T_28024 = _T_28021 & _T_28023; // @[LoadQueue.scala 327:31:@11692.4]
  assign _T_28025 = _T_28024 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@11693.4]
  assign _T_28026 = outputPriorityPorts_1_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@11694.4]
  assign _T_28029 = _T_28026 & _T_28023; // @[LoadQueue.scala 327:31:@11696.4]
  assign _T_28030 = _T_28029 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@11697.4]
  assign loadCompleting_2 = _T_28025 | _T_28030; // @[LoadQueue.scala 328:51:@11702.4]
  assign _T_28042 = outputPriorityPorts_0_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@11704.4]
  assign _T_28044 = loadCompleted_3 == 1'h0; // @[LoadQueue.scala 327:34:@11705.4]
  assign _T_28045 = _T_28042 & _T_28044; // @[LoadQueue.scala 327:31:@11706.4]
  assign _T_28046 = _T_28045 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@11707.4]
  assign _T_28047 = outputPriorityPorts_1_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@11708.4]
  assign _T_28050 = _T_28047 & _T_28044; // @[LoadQueue.scala 327:31:@11710.4]
  assign _T_28051 = _T_28050 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@11711.4]
  assign loadCompleting_3 = _T_28046 | _T_28051; // @[LoadQueue.scala 328:51:@11716.4]
  assign _T_28063 = outputPriorityPorts_0_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@11718.4]
  assign _T_28065 = loadCompleted_4 == 1'h0; // @[LoadQueue.scala 327:34:@11719.4]
  assign _T_28066 = _T_28063 & _T_28065; // @[LoadQueue.scala 327:31:@11720.4]
  assign _T_28067 = _T_28066 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@11721.4]
  assign _T_28068 = outputPriorityPorts_1_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@11722.4]
  assign _T_28071 = _T_28068 & _T_28065; // @[LoadQueue.scala 327:31:@11724.4]
  assign _T_28072 = _T_28071 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@11725.4]
  assign loadCompleting_4 = _T_28067 | _T_28072; // @[LoadQueue.scala 328:51:@11730.4]
  assign _T_28084 = outputPriorityPorts_0_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@11732.4]
  assign _T_28086 = loadCompleted_5 == 1'h0; // @[LoadQueue.scala 327:34:@11733.4]
  assign _T_28087 = _T_28084 & _T_28086; // @[LoadQueue.scala 327:31:@11734.4]
  assign _T_28088 = _T_28087 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@11735.4]
  assign _T_28089 = outputPriorityPorts_1_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@11736.4]
  assign _T_28092 = _T_28089 & _T_28086; // @[LoadQueue.scala 327:31:@11738.4]
  assign _T_28093 = _T_28092 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@11739.4]
  assign loadCompleting_5 = _T_28088 | _T_28093; // @[LoadQueue.scala 328:51:@11744.4]
  assign _T_28105 = outputPriorityPorts_0_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@11746.4]
  assign _T_28107 = loadCompleted_6 == 1'h0; // @[LoadQueue.scala 327:34:@11747.4]
  assign _T_28108 = _T_28105 & _T_28107; // @[LoadQueue.scala 327:31:@11748.4]
  assign _T_28109 = _T_28108 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@11749.4]
  assign _T_28110 = outputPriorityPorts_1_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@11750.4]
  assign _T_28113 = _T_28110 & _T_28107; // @[LoadQueue.scala 327:31:@11752.4]
  assign _T_28114 = _T_28113 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@11753.4]
  assign loadCompleting_6 = _T_28109 | _T_28114; // @[LoadQueue.scala 328:51:@11758.4]
  assign _T_28126 = outputPriorityPorts_0_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@11760.4]
  assign _T_28128 = loadCompleted_7 == 1'h0; // @[LoadQueue.scala 327:34:@11761.4]
  assign _T_28129 = _T_28126 & _T_28128; // @[LoadQueue.scala 327:31:@11762.4]
  assign _T_28130 = _T_28129 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@11763.4]
  assign _T_28131 = outputPriorityPorts_1_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@11764.4]
  assign _T_28134 = _T_28131 & _T_28128; // @[LoadQueue.scala 327:31:@11766.4]
  assign _T_28135 = _T_28134 & io_loadPorts_1_ready; // @[LoadQueue.scala 327:63:@11767.4]
  assign loadCompleting_7 = _T_28130 | _T_28135; // @[LoadQueue.scala 328:51:@11772.4]
  assign _GEN_658 = loadCompleting_0 ? 1'h1 : loadCompleted_0; // @[LoadQueue.scala 337:46:@11778.6]
  assign _GEN_659 = initBits_0 ? 1'h0 : _GEN_658; // @[LoadQueue.scala 335:34:@11774.4]
  assign _GEN_660 = loadCompleting_1 ? 1'h1 : loadCompleted_1; // @[LoadQueue.scala 337:46:@11785.6]
  assign _GEN_661 = initBits_1 ? 1'h0 : _GEN_660; // @[LoadQueue.scala 335:34:@11781.4]
  assign _GEN_662 = loadCompleting_2 ? 1'h1 : loadCompleted_2; // @[LoadQueue.scala 337:46:@11792.6]
  assign _GEN_663 = initBits_2 ? 1'h0 : _GEN_662; // @[LoadQueue.scala 335:34:@11788.4]
  assign _GEN_664 = loadCompleting_3 ? 1'h1 : loadCompleted_3; // @[LoadQueue.scala 337:46:@11799.6]
  assign _GEN_665 = initBits_3 ? 1'h0 : _GEN_664; // @[LoadQueue.scala 335:34:@11795.4]
  assign _GEN_666 = loadCompleting_4 ? 1'h1 : loadCompleted_4; // @[LoadQueue.scala 337:46:@11806.6]
  assign _GEN_667 = initBits_4 ? 1'h0 : _GEN_666; // @[LoadQueue.scala 335:34:@11802.4]
  assign _GEN_668 = loadCompleting_5 ? 1'h1 : loadCompleted_5; // @[LoadQueue.scala 337:46:@11813.6]
  assign _GEN_669 = initBits_5 ? 1'h0 : _GEN_668; // @[LoadQueue.scala 335:34:@11809.4]
  assign _GEN_670 = loadCompleting_6 ? 1'h1 : loadCompleted_6; // @[LoadQueue.scala 337:46:@11820.6]
  assign _GEN_671 = initBits_6 ? 1'h0 : _GEN_670; // @[LoadQueue.scala 335:34:@11816.4]
  assign _GEN_672 = loadCompleting_7 ? 1'h1 : loadCompleted_7; // @[LoadQueue.scala 337:46:@11827.6]
  assign _GEN_673 = initBits_7 ? 1'h0 : _GEN_672; // @[LoadQueue.scala 335:34:@11823.4]
  assign _T_28211 = _T_27982 | _T_28003; // @[LoadQueue.scala 348:24:@11864.4]
  assign _T_28212 = _T_28211 | _T_28024; // @[LoadQueue.scala 348:24:@11865.4]
  assign _T_28213 = _T_28212 | _T_28045; // @[LoadQueue.scala 348:24:@11866.4]
  assign _T_28214 = _T_28213 | _T_28066; // @[LoadQueue.scala 348:24:@11867.4]
  assign _T_28215 = _T_28214 | _T_28087; // @[LoadQueue.scala 348:24:@11868.4]
  assign _T_28216 = _T_28215 | _T_28108; // @[LoadQueue.scala 348:24:@11869.4]
  assign _T_28217 = _T_28216 | _T_28129; // @[LoadQueue.scala 348:24:@11870.4]
  assign _T_28226 = _T_28108 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@11872.6]
  assign _T_28227 = _T_28087 ? 3'h5 : _T_28226; // @[Mux.scala 31:69:@11873.6]
  assign _T_28228 = _T_28066 ? 3'h4 : _T_28227; // @[Mux.scala 31:69:@11874.6]
  assign _T_28229 = _T_28045 ? 3'h3 : _T_28228; // @[Mux.scala 31:69:@11875.6]
  assign _T_28230 = _T_28024 ? 3'h2 : _T_28229; // @[Mux.scala 31:69:@11876.6]
  assign _T_28231 = _T_28003 ? 3'h1 : _T_28230; // @[Mux.scala 31:69:@11877.6]
  assign _T_28232 = _T_27982 ? 3'h0 : _T_28231; // @[Mux.scala 31:69:@11878.6]
  assign _GEN_675 = 3'h1 == _T_28232 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@11879.6]
  assign _GEN_676 = 3'h2 == _T_28232 ? dataQ_2 : _GEN_675; // @[LoadQueue.scala 349:37:@11879.6]
  assign _GEN_677 = 3'h3 == _T_28232 ? dataQ_3 : _GEN_676; // @[LoadQueue.scala 349:37:@11879.6]
  assign _GEN_678 = 3'h4 == _T_28232 ? dataQ_4 : _GEN_677; // @[LoadQueue.scala 349:37:@11879.6]
  assign _GEN_679 = 3'h5 == _T_28232 ? dataQ_5 : _GEN_678; // @[LoadQueue.scala 349:37:@11879.6]
  assign _GEN_680 = 3'h6 == _T_28232 ? dataQ_6 : _GEN_679; // @[LoadQueue.scala 349:37:@11879.6]
  assign _GEN_681 = 3'h7 == _T_28232 ? dataQ_7 : _GEN_680; // @[LoadQueue.scala 349:37:@11879.6]
  assign _T_28287 = _T_27987 | _T_28008; // @[LoadQueue.scala 348:24:@11920.4]
  assign _T_28288 = _T_28287 | _T_28029; // @[LoadQueue.scala 348:24:@11921.4]
  assign _T_28289 = _T_28288 | _T_28050; // @[LoadQueue.scala 348:24:@11922.4]
  assign _T_28290 = _T_28289 | _T_28071; // @[LoadQueue.scala 348:24:@11923.4]
  assign _T_28291 = _T_28290 | _T_28092; // @[LoadQueue.scala 348:24:@11924.4]
  assign _T_28292 = _T_28291 | _T_28113; // @[LoadQueue.scala 348:24:@11925.4]
  assign _T_28293 = _T_28292 | _T_28134; // @[LoadQueue.scala 348:24:@11926.4]
  assign _T_28302 = _T_28113 ? 3'h6 : 3'h7; // @[Mux.scala 31:69:@11928.6]
  assign _T_28303 = _T_28092 ? 3'h5 : _T_28302; // @[Mux.scala 31:69:@11929.6]
  assign _T_28304 = _T_28071 ? 3'h4 : _T_28303; // @[Mux.scala 31:69:@11930.6]
  assign _T_28305 = _T_28050 ? 3'h3 : _T_28304; // @[Mux.scala 31:69:@11931.6]
  assign _T_28306 = _T_28029 ? 3'h2 : _T_28305; // @[Mux.scala 31:69:@11932.6]
  assign _T_28307 = _T_28008 ? 3'h1 : _T_28306; // @[Mux.scala 31:69:@11933.6]
  assign _T_28308 = _T_27987 ? 3'h0 : _T_28307; // @[Mux.scala 31:69:@11934.6]
  assign _GEN_685 = 3'h1 == _T_28308 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@11935.6]
  assign _GEN_686 = 3'h2 == _T_28308 ? dataQ_2 : _GEN_685; // @[LoadQueue.scala 349:37:@11935.6]
  assign _GEN_687 = 3'h3 == _T_28308 ? dataQ_3 : _GEN_686; // @[LoadQueue.scala 349:37:@11935.6]
  assign _GEN_688 = 3'h4 == _T_28308 ? dataQ_4 : _GEN_687; // @[LoadQueue.scala 349:37:@11935.6]
  assign _GEN_689 = 3'h5 == _T_28308 ? dataQ_5 : _GEN_688; // @[LoadQueue.scala 349:37:@11935.6]
  assign _GEN_690 = 3'h6 == _T_28308 ? dataQ_6 : _GEN_689; // @[LoadQueue.scala 349:37:@11935.6]
  assign _GEN_691 = 3'h7 == _T_28308 ? dataQ_7 : _GEN_690; // @[LoadQueue.scala 349:37:@11935.6]
  assign _GEN_695 = 3'h1 == head ? loadCompleted_1 : loadCompleted_0; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_696 = 3'h2 == head ? loadCompleted_2 : _GEN_695; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_697 = 3'h3 == head ? loadCompleted_3 : _GEN_696; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_698 = 3'h4 == head ? loadCompleted_4 : _GEN_697; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_699 = 3'h5 == head ? loadCompleted_5 : _GEN_698; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_700 = 3'h6 == head ? loadCompleted_6 : _GEN_699; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_701 = 3'h7 == head ? loadCompleted_7 : _GEN_700; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_703 = 3'h1 == head ? loadCompleting_1 : loadCompleting_0; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_704 = 3'h2 == head ? loadCompleting_2 : _GEN_703; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_705 = 3'h3 == head ? loadCompleting_3 : _GEN_704; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_706 = 3'h4 == head ? loadCompleting_4 : _GEN_705; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_707 = 3'h5 == head ? loadCompleting_5 : _GEN_706; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_708 = 3'h6 == head ? loadCompleting_6 : _GEN_707; // @[LoadQueue.scala 363:29:@11942.4]
  assign _GEN_709 = 3'h7 == head ? loadCompleting_7 : _GEN_708; // @[LoadQueue.scala 363:29:@11942.4]
  assign _T_28319 = _GEN_701 | _GEN_709; // @[LoadQueue.scala 363:29:@11942.4]
  assign _T_28320 = head != tail; // @[LoadQueue.scala 363:63:@11943.4]
  assign _T_28322 = io_loadEmpty == 1'h0; // @[LoadQueue.scala 363:75:@11944.4]
  assign _T_28323 = _T_28320 | _T_28322; // @[LoadQueue.scala 363:72:@11945.4]
  assign _T_28324 = _T_28319 & _T_28323; // @[LoadQueue.scala 363:54:@11946.4]
  assign _T_28327 = head + 3'h1; // @[util.scala 10:8:@11948.6]
  assign _GEN_144 = _T_28327 % 4'h8; // @[util.scala 10:14:@11949.6]
  assign _T_28328 = _GEN_144[3:0]; // @[util.scala 10:14:@11949.6]
  assign _GEN_710 = _T_28324 ? _T_28328 : {{1'd0}, head}; // @[LoadQueue.scala 363:91:@11947.4]
  assign _GEN_760 = {{1'd0}, io_bbNumLoads}; // @[util.scala 10:8:@11953.6]
  assign _T_28330 = tail + _GEN_760; // @[util.scala 10:8:@11953.6]
  assign _GEN_145 = _T_28330 % 4'h8; // @[util.scala 10:14:@11954.6]
  assign _T_28331 = _GEN_145[3:0]; // @[util.scala 10:14:@11954.6]
  assign _GEN_711 = io_bbStart ? _T_28331 : {{1'd0}, tail}; // @[LoadQueue.scala 367:20:@11952.4]
  assign _T_28333 = allocatedEntries_0 == 1'h0; // @[LoadQueue.scala 371:82:@11957.4]
  assign _T_28334 = loadCompleted_0 | _T_28333; // @[LoadQueue.scala 371:79:@11958.4]
  assign _T_28336 = allocatedEntries_1 == 1'h0; // @[LoadQueue.scala 371:82:@11959.4]
  assign _T_28337 = loadCompleted_1 | _T_28336; // @[LoadQueue.scala 371:79:@11960.4]
  assign _T_28339 = allocatedEntries_2 == 1'h0; // @[LoadQueue.scala 371:82:@11961.4]
  assign _T_28340 = loadCompleted_2 | _T_28339; // @[LoadQueue.scala 371:79:@11962.4]
  assign _T_28342 = allocatedEntries_3 == 1'h0; // @[LoadQueue.scala 371:82:@11963.4]
  assign _T_28343 = loadCompleted_3 | _T_28342; // @[LoadQueue.scala 371:79:@11964.4]
  assign _T_28345 = allocatedEntries_4 == 1'h0; // @[LoadQueue.scala 371:82:@11965.4]
  assign _T_28346 = loadCompleted_4 | _T_28345; // @[LoadQueue.scala 371:79:@11966.4]
  assign _T_28348 = allocatedEntries_5 == 1'h0; // @[LoadQueue.scala 371:82:@11967.4]
  assign _T_28349 = loadCompleted_5 | _T_28348; // @[LoadQueue.scala 371:79:@11968.4]
  assign _T_28351 = allocatedEntries_6 == 1'h0; // @[LoadQueue.scala 371:82:@11969.4]
  assign _T_28352 = loadCompleted_6 | _T_28351; // @[LoadQueue.scala 371:79:@11970.4]
  assign _T_28354 = allocatedEntries_7 == 1'h0; // @[LoadQueue.scala 371:82:@11971.4]
  assign _T_28355 = loadCompleted_7 | _T_28354; // @[LoadQueue.scala 371:79:@11972.4]
  assign _T_28372 = _T_28334 & _T_28337; // @[LoadQueue.scala 371:96:@11983.4]
  assign _T_28373 = _T_28372 & _T_28340; // @[LoadQueue.scala 371:96:@11984.4]
  assign _T_28374 = _T_28373 & _T_28343; // @[LoadQueue.scala 371:96:@11985.4]
  assign _T_28375 = _T_28374 & _T_28346; // @[LoadQueue.scala 371:96:@11986.4]
  assign _T_28376 = _T_28375 & _T_28349; // @[LoadQueue.scala 371:96:@11987.4]
  assign _T_28377 = _T_28376 & _T_28352; // @[LoadQueue.scala 371:96:@11988.4]
  assign io_loadTail = tail; // @[LoadQueue.scala 380:15:@11992.4]
  assign io_loadHead = head; // @[LoadQueue.scala 379:15:@11991.4]
  assign io_loadEmpty = _T_28377 & _T_28355; // @[LoadQueue.scala 371:16:@11990.4]
  assign io_loadAddrDone_0 = addrKnown_0; // @[LoadQueue.scala 382:19:@12001.4]
  assign io_loadAddrDone_1 = addrKnown_1; // @[LoadQueue.scala 382:19:@12002.4]
  assign io_loadAddrDone_2 = addrKnown_2; // @[LoadQueue.scala 382:19:@12003.4]
  assign io_loadAddrDone_3 = addrKnown_3; // @[LoadQueue.scala 382:19:@12004.4]
  assign io_loadAddrDone_4 = addrKnown_4; // @[LoadQueue.scala 382:19:@12005.4]
  assign io_loadAddrDone_5 = addrKnown_5; // @[LoadQueue.scala 382:19:@12006.4]
  assign io_loadAddrDone_6 = addrKnown_6; // @[LoadQueue.scala 382:19:@12007.4]
  assign io_loadAddrDone_7 = addrKnown_7; // @[LoadQueue.scala 382:19:@12008.4]
  assign io_loadDataDone_0 = dataKnown_0; // @[LoadQueue.scala 383:19:@12009.4]
  assign io_loadDataDone_1 = dataKnown_1; // @[LoadQueue.scala 383:19:@12010.4]
  assign io_loadDataDone_2 = dataKnown_2; // @[LoadQueue.scala 383:19:@12011.4]
  assign io_loadDataDone_3 = dataKnown_3; // @[LoadQueue.scala 383:19:@12012.4]
  assign io_loadDataDone_4 = dataKnown_4; // @[LoadQueue.scala 383:19:@12013.4]
  assign io_loadDataDone_5 = dataKnown_5; // @[LoadQueue.scala 383:19:@12014.4]
  assign io_loadDataDone_6 = dataKnown_6; // @[LoadQueue.scala 383:19:@12015.4]
  assign io_loadDataDone_7 = dataKnown_7; // @[LoadQueue.scala 383:19:@12016.4]
  assign io_loadAddrQueue_0 = addrQ_0; // @[LoadQueue.scala 381:20:@11993.4]
  assign io_loadAddrQueue_1 = addrQ_1; // @[LoadQueue.scala 381:20:@11994.4]
  assign io_loadAddrQueue_2 = addrQ_2; // @[LoadQueue.scala 381:20:@11995.4]
  assign io_loadAddrQueue_3 = addrQ_3; // @[LoadQueue.scala 381:20:@11996.4]
  assign io_loadAddrQueue_4 = addrQ_4; // @[LoadQueue.scala 381:20:@11997.4]
  assign io_loadAddrQueue_5 = addrQ_5; // @[LoadQueue.scala 381:20:@11998.4]
  assign io_loadAddrQueue_6 = addrQ_6; // @[LoadQueue.scala 381:20:@11999.4]
  assign io_loadAddrQueue_7 = addrQ_7; // @[LoadQueue.scala 381:20:@12000.4]
  assign io_loadPorts_0_valid = _T_28216 | _T_28129; // @[LoadQueue.scala 350:38:@11880.6 LoadQueue.scala 353:38:@11884.6]
  assign io_loadPorts_0_bits = _T_28217 ? _GEN_681 : 32'h0; // @[LoadQueue.scala 349:37:@11879.6 LoadQueue.scala 352:37:@11883.6]
  assign io_loadPorts_1_valid = _T_28292 | _T_28134; // @[LoadQueue.scala 350:38:@11936.6 LoadQueue.scala 353:38:@11940.6]
  assign io_loadPorts_1_bits = _T_28293 ? _GEN_691 : 32'h0; // @[LoadQueue.scala 349:37:@11935.6 LoadQueue.scala 352:37:@11939.6]
  assign io_loadAddrToMem = _T_25202 ? _GEN_575 : 32'h0; // @[LoadQueue.scala 248:24:@10033.6 LoadQueue.scala 251:24:@10037.6]
  assign io_loadEnableToMem = _T_25201 | loadRequest_7; // @[LoadQueue.scala 246:22:@10016.4 LoadQueue.scala 249:26:@10034.6 LoadQueue.scala 252:26:@10038.6]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  portQ_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  portQ_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  portQ_2 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  portQ_3 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  portQ_4 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  portQ_5 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  portQ_6 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  portQ_7 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  addrQ_0 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  addrQ_1 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  addrQ_2 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  addrQ_3 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  addrQ_4 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  addrQ_5 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  addrQ_6 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  addrQ_7 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  dataQ_0 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  dataQ_1 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  dataQ_2 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  dataQ_3 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  dataQ_4 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  dataQ_5 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  dataQ_6 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  dataQ_7 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrKnown_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrKnown_1 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrKnown_2 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrKnown_3 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrKnown_4 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrKnown_5 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrKnown_6 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrKnown_7 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  dataKnown_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  dataKnown_1 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  dataKnown_2 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  dataKnown_3 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  dataKnown_4 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  dataKnown_5 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  dataKnown_6 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  dataKnown_7 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  loadCompleted_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  loadCompleted_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  loadCompleted_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  loadCompleted_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  loadCompleted_4 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  loadCompleted_5 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  loadCompleted_6 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  loadCompleted_7 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  bypassInitiated_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  bypassInitiated_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  bypassInitiated_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  bypassInitiated_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  bypassInitiated_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  bypassInitiated_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  bypassInitiated_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  bypassInitiated_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  checkBits_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  checkBits_1 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  checkBits_2 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  checkBits_3 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  checkBits_4 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  checkBits_5 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  checkBits_6 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  checkBits_7 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  previousStoreHead = _RAND_82[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  conflictPReg_0_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  conflictPReg_0_1 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  conflictPReg_0_2 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  conflictPReg_0_3 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  conflictPReg_0_4 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  conflictPReg_0_5 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  conflictPReg_0_6 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  conflictPReg_0_7 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  conflictPReg_1_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  conflictPReg_1_1 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  conflictPReg_1_2 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  conflictPReg_1_3 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  conflictPReg_1_4 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  conflictPReg_1_5 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  conflictPReg_1_6 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  conflictPReg_1_7 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  conflictPReg_2_0 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  conflictPReg_2_1 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  conflictPReg_2_2 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  conflictPReg_2_3 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  conflictPReg_2_4 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  conflictPReg_2_5 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  conflictPReg_2_6 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  conflictPReg_2_7 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  conflictPReg_3_0 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  conflictPReg_3_1 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  conflictPReg_3_2 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  conflictPReg_3_3 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  conflictPReg_3_4 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  conflictPReg_3_5 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  conflictPReg_3_6 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  conflictPReg_3_7 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  conflictPReg_4_0 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  conflictPReg_4_1 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  conflictPReg_4_2 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  conflictPReg_4_3 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  conflictPReg_4_4 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  conflictPReg_4_5 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  conflictPReg_4_6 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  conflictPReg_4_7 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  conflictPReg_5_0 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  conflictPReg_5_1 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  conflictPReg_5_2 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  conflictPReg_5_3 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  conflictPReg_5_4 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  conflictPReg_5_5 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  conflictPReg_5_6 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  conflictPReg_5_7 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  conflictPReg_6_0 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  conflictPReg_6_1 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  conflictPReg_6_2 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  conflictPReg_6_3 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  conflictPReg_6_4 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  conflictPReg_6_5 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  conflictPReg_6_6 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  conflictPReg_6_7 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  conflictPReg_7_0 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  conflictPReg_7_1 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  conflictPReg_7_2 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  conflictPReg_7_3 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  conflictPReg_7_4 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  conflictPReg_7_5 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  conflictPReg_7_6 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  conflictPReg_7_7 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_0 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_1 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_2 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_3 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_4 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_5 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_6 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_7 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_0 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_1 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_2 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_3 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_4 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_5 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_6 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_7 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_0 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_1 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_2 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_3 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_4 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_5 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_6 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_7 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_0 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_1 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_2 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_3 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_4 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_5 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_6 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_7 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_0 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_1 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_2 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_3 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_4 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_5 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_6 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_7 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_0 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_1 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_2 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_3 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_4 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_5 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_6 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_7 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_0 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_1 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_2 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_3 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_4 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_5 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_6 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_7 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_0 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_1 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_2 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_3 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_4 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_5 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_6 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_7 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_0 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_1 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_2 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_3 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_4 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_5 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_6 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_7 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  shiftedStoreDataQPreg_0 = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  shiftedStoreDataQPreg_1 = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  shiftedStoreDataQPreg_2 = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  shiftedStoreDataQPreg_3 = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  shiftedStoreDataQPreg_4 = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  shiftedStoreDataQPreg_5 = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  shiftedStoreDataQPreg_6 = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  shiftedStoreDataQPreg_7 = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  addrKnownPReg_0 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  addrKnownPReg_1 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  addrKnownPReg_2 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  addrKnownPReg_3 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  addrKnownPReg_4 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  addrKnownPReg_5 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  addrKnownPReg_6 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  addrKnownPReg_7 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  dataKnownPReg_0 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  dataKnownPReg_1 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  dataKnownPReg_2 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  dataKnownPReg_3 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  dataKnownPReg_4 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  dataKnownPReg_5 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  dataKnownPReg_6 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  dataKnownPReg_7 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  prevPriorityRequest_7 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  prevPriorityRequest_6 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  prevPriorityRequest_5 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  prevPriorityRequest_4 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  prevPriorityRequest_3 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  prevPriorityRequest_2 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  prevPriorityRequest_1 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  prevPriorityRequest_0 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 3'h0;
    end else begin
      head <= _GEN_710[2:0];
    end
    if (reset) begin
      tail <= 3'h0;
    end else begin
      tail <= _GEN_711[2:0];
    end
    if (reset) begin
      offsetQ_0 <= 3'h0;
    end else begin
      if (initBits_0) begin
        if (3'h7 == _T_1132) begin
          offsetQ_0 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1132) begin
            offsetQ_0 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1132) begin
              offsetQ_0 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1132) begin
                offsetQ_0 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1132) begin
                  offsetQ_0 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1132) begin
                    offsetQ_0 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1132) begin
                      offsetQ_0 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_0 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 3'h0;
    end else begin
      if (initBits_1) begin
        if (3'h7 == _T_1150) begin
          offsetQ_1 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1150) begin
            offsetQ_1 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1150) begin
              offsetQ_1 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1150) begin
                offsetQ_1 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1150) begin
                  offsetQ_1 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1150) begin
                    offsetQ_1 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1150) begin
                      offsetQ_1 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_1 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 3'h0;
    end else begin
      if (initBits_2) begin
        if (3'h7 == _T_1168) begin
          offsetQ_2 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1168) begin
            offsetQ_2 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1168) begin
              offsetQ_2 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1168) begin
                offsetQ_2 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1168) begin
                  offsetQ_2 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1168) begin
                    offsetQ_2 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1168) begin
                      offsetQ_2 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_2 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 3'h0;
    end else begin
      if (initBits_3) begin
        if (3'h7 == _T_1186) begin
          offsetQ_3 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1186) begin
            offsetQ_3 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1186) begin
              offsetQ_3 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1186) begin
                offsetQ_3 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1186) begin
                  offsetQ_3 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1186) begin
                    offsetQ_3 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1186) begin
                      offsetQ_3 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_3 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 3'h0;
    end else begin
      if (initBits_4) begin
        if (3'h7 == _T_1204) begin
          offsetQ_4 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1204) begin
            offsetQ_4 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1204) begin
              offsetQ_4 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1204) begin
                offsetQ_4 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1204) begin
                  offsetQ_4 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1204) begin
                    offsetQ_4 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1204) begin
                      offsetQ_4 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_4 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 3'h0;
    end else begin
      if (initBits_5) begin
        if (3'h7 == _T_1222) begin
          offsetQ_5 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1222) begin
            offsetQ_5 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1222) begin
              offsetQ_5 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1222) begin
                offsetQ_5 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1222) begin
                  offsetQ_5 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1222) begin
                    offsetQ_5 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1222) begin
                      offsetQ_5 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_5 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 3'h0;
    end else begin
      if (initBits_6) begin
        if (3'h7 == _T_1240) begin
          offsetQ_6 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1240) begin
            offsetQ_6 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1240) begin
              offsetQ_6 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1240) begin
                offsetQ_6 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1240) begin
                  offsetQ_6 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1240) begin
                    offsetQ_6 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1240) begin
                      offsetQ_6 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_6 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 3'h0;
    end else begin
      if (initBits_7) begin
        if (3'h7 == _T_1258) begin
          offsetQ_7 <= io_bbLoadOffsets_7;
        end else begin
          if (3'h6 == _T_1258) begin
            offsetQ_7 <= io_bbLoadOffsets_6;
          end else begin
            if (3'h5 == _T_1258) begin
              offsetQ_7 <= io_bbLoadOffsets_5;
            end else begin
              if (3'h4 == _T_1258) begin
                offsetQ_7 <= io_bbLoadOffsets_4;
              end else begin
                if (3'h3 == _T_1258) begin
                  offsetQ_7 <= io_bbLoadOffsets_3;
                end else begin
                  if (3'h2 == _T_1258) begin
                    offsetQ_7 <= io_bbLoadOffsets_2;
                  end else begin
                    if (3'h1 == _T_1258) begin
                      offsetQ_7 <= io_bbLoadOffsets_1;
                    end else begin
                      offsetQ_7 <= io_bbLoadOffsets_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        if (3'h7 == _T_1132) begin
          portQ_0 <= 1'h0;
        end else begin
          if (3'h6 == _T_1132) begin
            portQ_0 <= 1'h0;
          end else begin
            if (3'h5 == _T_1132) begin
              portQ_0 <= 1'h0;
            end else begin
              if (3'h4 == _T_1132) begin
                portQ_0 <= 1'h0;
              end else begin
                if (3'h3 == _T_1132) begin
                  portQ_0 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1132) begin
                    portQ_0 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1132) begin
                      portQ_0 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_0 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        if (3'h7 == _T_1150) begin
          portQ_1 <= 1'h0;
        end else begin
          if (3'h6 == _T_1150) begin
            portQ_1 <= 1'h0;
          end else begin
            if (3'h5 == _T_1150) begin
              portQ_1 <= 1'h0;
            end else begin
              if (3'h4 == _T_1150) begin
                portQ_1 <= 1'h0;
              end else begin
                if (3'h3 == _T_1150) begin
                  portQ_1 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1150) begin
                    portQ_1 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1150) begin
                      portQ_1 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_1 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        if (3'h7 == _T_1168) begin
          portQ_2 <= 1'h0;
        end else begin
          if (3'h6 == _T_1168) begin
            portQ_2 <= 1'h0;
          end else begin
            if (3'h5 == _T_1168) begin
              portQ_2 <= 1'h0;
            end else begin
              if (3'h4 == _T_1168) begin
                portQ_2 <= 1'h0;
              end else begin
                if (3'h3 == _T_1168) begin
                  portQ_2 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1168) begin
                    portQ_2 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1168) begin
                      portQ_2 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_2 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        if (3'h7 == _T_1186) begin
          portQ_3 <= 1'h0;
        end else begin
          if (3'h6 == _T_1186) begin
            portQ_3 <= 1'h0;
          end else begin
            if (3'h5 == _T_1186) begin
              portQ_3 <= 1'h0;
            end else begin
              if (3'h4 == _T_1186) begin
                portQ_3 <= 1'h0;
              end else begin
                if (3'h3 == _T_1186) begin
                  portQ_3 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1186) begin
                    portQ_3 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1186) begin
                      portQ_3 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_3 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        if (3'h7 == _T_1204) begin
          portQ_4 <= 1'h0;
        end else begin
          if (3'h6 == _T_1204) begin
            portQ_4 <= 1'h0;
          end else begin
            if (3'h5 == _T_1204) begin
              portQ_4 <= 1'h0;
            end else begin
              if (3'h4 == _T_1204) begin
                portQ_4 <= 1'h0;
              end else begin
                if (3'h3 == _T_1204) begin
                  portQ_4 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1204) begin
                    portQ_4 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1204) begin
                      portQ_4 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_4 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        if (3'h7 == _T_1222) begin
          portQ_5 <= 1'h0;
        end else begin
          if (3'h6 == _T_1222) begin
            portQ_5 <= 1'h0;
          end else begin
            if (3'h5 == _T_1222) begin
              portQ_5 <= 1'h0;
            end else begin
              if (3'h4 == _T_1222) begin
                portQ_5 <= 1'h0;
              end else begin
                if (3'h3 == _T_1222) begin
                  portQ_5 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1222) begin
                    portQ_5 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1222) begin
                      portQ_5 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_5 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        if (3'h7 == _T_1240) begin
          portQ_6 <= 1'h0;
        end else begin
          if (3'h6 == _T_1240) begin
            portQ_6 <= 1'h0;
          end else begin
            if (3'h5 == _T_1240) begin
              portQ_6 <= 1'h0;
            end else begin
              if (3'h4 == _T_1240) begin
                portQ_6 <= 1'h0;
              end else begin
                if (3'h3 == _T_1240) begin
                  portQ_6 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1240) begin
                    portQ_6 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1240) begin
                      portQ_6 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_6 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        if (3'h7 == _T_1258) begin
          portQ_7 <= 1'h0;
        end else begin
          if (3'h6 == _T_1258) begin
            portQ_7 <= 1'h0;
          end else begin
            if (3'h5 == _T_1258) begin
              portQ_7 <= 1'h0;
            end else begin
              if (3'h4 == _T_1258) begin
                portQ_7 <= 1'h0;
              end else begin
                if (3'h3 == _T_1258) begin
                  portQ_7 <= 1'h0;
                end else begin
                  if (3'h2 == _T_1258) begin
                    portQ_7 <= 1'h0;
                  end else begin
                    if (3'h1 == _T_1258) begin
                      portQ_7 <= io_bbLoadPorts_1;
                    end else begin
                      portQ_7 <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_27835) begin
          if (_T_27837) begin
            addrQ_0 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_0 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_27853) begin
          if (_T_27855) begin
            addrQ_1 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_1 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_27871) begin
          if (_T_27873) begin
            addrQ_2 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_2 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_27889) begin
          if (_T_27891) begin
            addrQ_3 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_3 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_27907) begin
          if (_T_27909) begin
            addrQ_4 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_4 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_27925) begin
          if (_T_27927) begin
            addrQ_5 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_5 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_27943) begin
          if (_T_27945) begin
            addrQ_6 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_6 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_27961) begin
          if (_T_27963) begin
            addrQ_7 <= io_addrFromLoadPorts_1;
          end else begin
            addrQ_7 <= io_addrFromLoadPorts_0;
          end
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (bypassRequest_0) begin
        if (_T_23546) begin
          if (3'h7 == _T_23537) begin
            dataQ_0 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23537) begin
              dataQ_0 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23537) begin
                dataQ_0 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23537) begin
                  dataQ_0 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23537) begin
                    dataQ_0 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23537) begin
                      dataQ_0 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23537) begin
                        dataQ_0 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_0 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_0 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_0) begin
          dataQ_0 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (bypassRequest_1) begin
        if (_T_23626) begin
          if (3'h7 == _T_23617) begin
            dataQ_1 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23617) begin
              dataQ_1 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23617) begin
                dataQ_1 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23617) begin
                  dataQ_1 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23617) begin
                    dataQ_1 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23617) begin
                      dataQ_1 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23617) begin
                        dataQ_1 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_1 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_1 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_1) begin
          dataQ_1 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (bypassRequest_2) begin
        if (_T_23706) begin
          if (3'h7 == _T_23697) begin
            dataQ_2 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23697) begin
              dataQ_2 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23697) begin
                dataQ_2 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23697) begin
                  dataQ_2 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23697) begin
                    dataQ_2 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23697) begin
                      dataQ_2 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23697) begin
                        dataQ_2 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_2 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_2 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_2) begin
          dataQ_2 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (bypassRequest_3) begin
        if (_T_23786) begin
          if (3'h7 == _T_23777) begin
            dataQ_3 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23777) begin
              dataQ_3 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23777) begin
                dataQ_3 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23777) begin
                  dataQ_3 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23777) begin
                    dataQ_3 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23777) begin
                      dataQ_3 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23777) begin
                        dataQ_3 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_3 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_3 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_3) begin
          dataQ_3 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (bypassRequest_4) begin
        if (_T_23866) begin
          if (3'h7 == _T_23857) begin
            dataQ_4 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23857) begin
              dataQ_4 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23857) begin
                dataQ_4 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23857) begin
                  dataQ_4 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23857) begin
                    dataQ_4 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23857) begin
                      dataQ_4 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23857) begin
                        dataQ_4 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_4 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_4 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_4) begin
          dataQ_4 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (bypassRequest_5) begin
        if (_T_23946) begin
          if (3'h7 == _T_23937) begin
            dataQ_5 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_23937) begin
              dataQ_5 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_23937) begin
                dataQ_5 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_23937) begin
                  dataQ_5 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_23937) begin
                    dataQ_5 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_23937) begin
                      dataQ_5 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_23937) begin
                        dataQ_5 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_5 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_5 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_5) begin
          dataQ_5 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (bypassRequest_6) begin
        if (_T_24026) begin
          if (3'h7 == _T_24017) begin
            dataQ_6 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_24017) begin
              dataQ_6 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_24017) begin
                dataQ_6 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_24017) begin
                  dataQ_6 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_24017) begin
                    dataQ_6 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_24017) begin
                      dataQ_6 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_24017) begin
                        dataQ_6 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_6 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_6 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_6) begin
          dataQ_6 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (bypassRequest_7) begin
        if (_T_24106) begin
          if (3'h7 == _T_24097) begin
            dataQ_7 <= shiftedStoreDataQPreg_7;
          end else begin
            if (3'h6 == _T_24097) begin
              dataQ_7 <= shiftedStoreDataQPreg_6;
            end else begin
              if (3'h5 == _T_24097) begin
                dataQ_7 <= shiftedStoreDataQPreg_5;
              end else begin
                if (3'h4 == _T_24097) begin
                  dataQ_7 <= shiftedStoreDataQPreg_4;
                end else begin
                  if (3'h3 == _T_24097) begin
                    dataQ_7 <= shiftedStoreDataQPreg_3;
                  end else begin
                    if (3'h2 == _T_24097) begin
                      dataQ_7 <= shiftedStoreDataQPreg_2;
                    end else begin
                      if (3'h1 == _T_24097) begin
                        dataQ_7 <= shiftedStoreDataQPreg_1;
                      end else begin
                        dataQ_7 <= shiftedStoreDataQPreg_0;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_7 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_7) begin
          dataQ_7 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_27835) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_27853) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_27871) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_27889) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_27907) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_27925) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_27943) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_27961) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_25225) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_25228) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_25231) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_25234) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_25237) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_25240) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_25243) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_25246) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        loadCompleted_0 <= 1'h0;
      end else begin
        if (loadCompleting_0) begin
          loadCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        loadCompleted_1 <= 1'h0;
      end else begin
        if (loadCompleting_1) begin
          loadCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        loadCompleted_2 <= 1'h0;
      end else begin
        if (loadCompleting_2) begin
          loadCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        loadCompleted_3 <= 1'h0;
      end else begin
        if (loadCompleting_3) begin
          loadCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        loadCompleted_4 <= 1'h0;
      end else begin
        if (loadCompleting_4) begin
          loadCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        loadCompleted_5 <= 1'h0;
      end else begin
        if (loadCompleting_5) begin
          loadCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        loadCompleted_6 <= 1'h0;
      end else begin
        if (loadCompleting_6) begin
          loadCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        loadCompleted_7 <= 1'h0;
      end else begin
        if (loadCompleting_7) begin
          loadCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1102;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1103;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1104;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1105;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1106;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1107;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1108;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1109;
    end
    if (reset) begin
      bypassInitiated_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        bypassInitiated_0 <= 1'h0;
      end else begin
        if (bypassRequest_0) begin
          bypassInitiated_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        bypassInitiated_1 <= 1'h0;
      end else begin
        if (bypassRequest_1) begin
          bypassInitiated_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        bypassInitiated_2 <= 1'h0;
      end else begin
        if (bypassRequest_2) begin
          bypassInitiated_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        bypassInitiated_3 <= 1'h0;
      end else begin
        if (bypassRequest_3) begin
          bypassInitiated_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        bypassInitiated_4 <= 1'h0;
      end else begin
        if (bypassRequest_4) begin
          bypassInitiated_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        bypassInitiated_5 <= 1'h0;
      end else begin
        if (bypassRequest_5) begin
          bypassInitiated_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        bypassInitiated_6 <= 1'h0;
      end else begin
        if (bypassRequest_6) begin
          bypassInitiated_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        bypassInitiated_7 <= 1'h0;
      end else begin
        if (bypassRequest_7) begin
          bypassInitiated_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_1285;
      end else begin
        if (io_storeEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_1289) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_1297) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_1315;
      end else begin
        if (io_storeEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_1319) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_1327) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_1345;
      end else begin
        if (io_storeEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_1349) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_1357) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_1375;
      end else begin
        if (io_storeEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_1379) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_1387) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_1405;
      end else begin
        if (io_storeEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_1409) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_1417) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_1435;
      end else begin
        if (io_storeEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_1439) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_1447) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_1465;
      end else begin
        if (io_storeEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_1469) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_1477) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_1495;
      end else begin
        if (io_storeEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_1499) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_1507) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    previousStoreHead <= io_storeHead;
    conflictPReg_0_0 <= _T_6194[0];
    conflictPReg_0_1 <= _T_6194[1];
    conflictPReg_0_2 <= _T_6194[2];
    conflictPReg_0_3 <= _T_6194[3];
    conflictPReg_0_4 <= _T_6194[4];
    conflictPReg_0_5 <= _T_6194[5];
    conflictPReg_0_6 <= _T_6194[6];
    conflictPReg_0_7 <= _T_6194[7];
    conflictPReg_1_0 <= _T_6508[0];
    conflictPReg_1_1 <= _T_6508[1];
    conflictPReg_1_2 <= _T_6508[2];
    conflictPReg_1_3 <= _T_6508[3];
    conflictPReg_1_4 <= _T_6508[4];
    conflictPReg_1_5 <= _T_6508[5];
    conflictPReg_1_6 <= _T_6508[6];
    conflictPReg_1_7 <= _T_6508[7];
    conflictPReg_2_0 <= _T_6822[0];
    conflictPReg_2_1 <= _T_6822[1];
    conflictPReg_2_2 <= _T_6822[2];
    conflictPReg_2_3 <= _T_6822[3];
    conflictPReg_2_4 <= _T_6822[4];
    conflictPReg_2_5 <= _T_6822[5];
    conflictPReg_2_6 <= _T_6822[6];
    conflictPReg_2_7 <= _T_6822[7];
    conflictPReg_3_0 <= _T_7136[0];
    conflictPReg_3_1 <= _T_7136[1];
    conflictPReg_3_2 <= _T_7136[2];
    conflictPReg_3_3 <= _T_7136[3];
    conflictPReg_3_4 <= _T_7136[4];
    conflictPReg_3_5 <= _T_7136[5];
    conflictPReg_3_6 <= _T_7136[6];
    conflictPReg_3_7 <= _T_7136[7];
    conflictPReg_4_0 <= _T_7450[0];
    conflictPReg_4_1 <= _T_7450[1];
    conflictPReg_4_2 <= _T_7450[2];
    conflictPReg_4_3 <= _T_7450[3];
    conflictPReg_4_4 <= _T_7450[4];
    conflictPReg_4_5 <= _T_7450[5];
    conflictPReg_4_6 <= _T_7450[6];
    conflictPReg_4_7 <= _T_7450[7];
    conflictPReg_5_0 <= _T_7764[0];
    conflictPReg_5_1 <= _T_7764[1];
    conflictPReg_5_2 <= _T_7764[2];
    conflictPReg_5_3 <= _T_7764[3];
    conflictPReg_5_4 <= _T_7764[4];
    conflictPReg_5_5 <= _T_7764[5];
    conflictPReg_5_6 <= _T_7764[6];
    conflictPReg_5_7 <= _T_7764[7];
    conflictPReg_6_0 <= _T_8078[0];
    conflictPReg_6_1 <= _T_8078[1];
    conflictPReg_6_2 <= _T_8078[2];
    conflictPReg_6_3 <= _T_8078[3];
    conflictPReg_6_4 <= _T_8078[4];
    conflictPReg_6_5 <= _T_8078[5];
    conflictPReg_6_6 <= _T_8078[6];
    conflictPReg_6_7 <= _T_8078[7];
    conflictPReg_7_0 <= _T_8392[0];
    conflictPReg_7_1 <= _T_8392[1];
    conflictPReg_7_2 <= _T_8392[2];
    conflictPReg_7_3 <= _T_8392[3];
    conflictPReg_7_4 <= _T_8392[4];
    conflictPReg_7_5 <= _T_8392[5];
    conflictPReg_7_6 <= _T_8392[6];
    conflictPReg_7_7 <= _T_8392[7];
    storeAddrNotKnownFlagsPReg_0_0 <= _T_14574[0];
    storeAddrNotKnownFlagsPReg_0_1 <= _T_14574[1];
    storeAddrNotKnownFlagsPReg_0_2 <= _T_14574[2];
    storeAddrNotKnownFlagsPReg_0_3 <= _T_14574[3];
    storeAddrNotKnownFlagsPReg_0_4 <= _T_14574[4];
    storeAddrNotKnownFlagsPReg_0_5 <= _T_14574[5];
    storeAddrNotKnownFlagsPReg_0_6 <= _T_14574[6];
    storeAddrNotKnownFlagsPReg_0_7 <= _T_14574[7];
    storeAddrNotKnownFlagsPReg_1_0 <= _T_14888[0];
    storeAddrNotKnownFlagsPReg_1_1 <= _T_14888[1];
    storeAddrNotKnownFlagsPReg_1_2 <= _T_14888[2];
    storeAddrNotKnownFlagsPReg_1_3 <= _T_14888[3];
    storeAddrNotKnownFlagsPReg_1_4 <= _T_14888[4];
    storeAddrNotKnownFlagsPReg_1_5 <= _T_14888[5];
    storeAddrNotKnownFlagsPReg_1_6 <= _T_14888[6];
    storeAddrNotKnownFlagsPReg_1_7 <= _T_14888[7];
    storeAddrNotKnownFlagsPReg_2_0 <= _T_15202[0];
    storeAddrNotKnownFlagsPReg_2_1 <= _T_15202[1];
    storeAddrNotKnownFlagsPReg_2_2 <= _T_15202[2];
    storeAddrNotKnownFlagsPReg_2_3 <= _T_15202[3];
    storeAddrNotKnownFlagsPReg_2_4 <= _T_15202[4];
    storeAddrNotKnownFlagsPReg_2_5 <= _T_15202[5];
    storeAddrNotKnownFlagsPReg_2_6 <= _T_15202[6];
    storeAddrNotKnownFlagsPReg_2_7 <= _T_15202[7];
    storeAddrNotKnownFlagsPReg_3_0 <= _T_15516[0];
    storeAddrNotKnownFlagsPReg_3_1 <= _T_15516[1];
    storeAddrNotKnownFlagsPReg_3_2 <= _T_15516[2];
    storeAddrNotKnownFlagsPReg_3_3 <= _T_15516[3];
    storeAddrNotKnownFlagsPReg_3_4 <= _T_15516[4];
    storeAddrNotKnownFlagsPReg_3_5 <= _T_15516[5];
    storeAddrNotKnownFlagsPReg_3_6 <= _T_15516[6];
    storeAddrNotKnownFlagsPReg_3_7 <= _T_15516[7];
    storeAddrNotKnownFlagsPReg_4_0 <= _T_15830[0];
    storeAddrNotKnownFlagsPReg_4_1 <= _T_15830[1];
    storeAddrNotKnownFlagsPReg_4_2 <= _T_15830[2];
    storeAddrNotKnownFlagsPReg_4_3 <= _T_15830[3];
    storeAddrNotKnownFlagsPReg_4_4 <= _T_15830[4];
    storeAddrNotKnownFlagsPReg_4_5 <= _T_15830[5];
    storeAddrNotKnownFlagsPReg_4_6 <= _T_15830[6];
    storeAddrNotKnownFlagsPReg_4_7 <= _T_15830[7];
    storeAddrNotKnownFlagsPReg_5_0 <= _T_16144[0];
    storeAddrNotKnownFlagsPReg_5_1 <= _T_16144[1];
    storeAddrNotKnownFlagsPReg_5_2 <= _T_16144[2];
    storeAddrNotKnownFlagsPReg_5_3 <= _T_16144[3];
    storeAddrNotKnownFlagsPReg_5_4 <= _T_16144[4];
    storeAddrNotKnownFlagsPReg_5_5 <= _T_16144[5];
    storeAddrNotKnownFlagsPReg_5_6 <= _T_16144[6];
    storeAddrNotKnownFlagsPReg_5_7 <= _T_16144[7];
    storeAddrNotKnownFlagsPReg_6_0 <= _T_16458[0];
    storeAddrNotKnownFlagsPReg_6_1 <= _T_16458[1];
    storeAddrNotKnownFlagsPReg_6_2 <= _T_16458[2];
    storeAddrNotKnownFlagsPReg_6_3 <= _T_16458[3];
    storeAddrNotKnownFlagsPReg_6_4 <= _T_16458[4];
    storeAddrNotKnownFlagsPReg_6_5 <= _T_16458[5];
    storeAddrNotKnownFlagsPReg_6_6 <= _T_16458[6];
    storeAddrNotKnownFlagsPReg_6_7 <= _T_16458[7];
    storeAddrNotKnownFlagsPReg_7_0 <= _T_16772[0];
    storeAddrNotKnownFlagsPReg_7_1 <= _T_16772[1];
    storeAddrNotKnownFlagsPReg_7_2 <= _T_16772[2];
    storeAddrNotKnownFlagsPReg_7_3 <= _T_16772[3];
    storeAddrNotKnownFlagsPReg_7_4 <= _T_16772[4];
    storeAddrNotKnownFlagsPReg_7_5 <= _T_16772[5];
    storeAddrNotKnownFlagsPReg_7_6 <= _T_16772[6];
    storeAddrNotKnownFlagsPReg_7_7 <= _T_16772[7];
    shiftedStoreDataKnownPReg_0 <= _T_2684[0];
    shiftedStoreDataKnownPReg_1 <= _T_2684[1];
    shiftedStoreDataKnownPReg_2 <= _T_2684[2];
    shiftedStoreDataKnownPReg_3 <= _T_2684[3];
    shiftedStoreDataKnownPReg_4 <= _T_2684[4];
    shiftedStoreDataKnownPReg_5 <= _T_2684[5];
    shiftedStoreDataKnownPReg_6 <= _T_2684[6];
    shiftedStoreDataKnownPReg_7 <= _T_2684[7];
    shiftedStoreDataQPreg_0 <= _T_2371[31:0];
    shiftedStoreDataQPreg_1 <= _T_2371[63:32];
    shiftedStoreDataQPreg_2 <= _T_2371[95:64];
    shiftedStoreDataQPreg_3 <= _T_2371[127:96];
    shiftedStoreDataQPreg_4 <= _T_2371[159:128];
    shiftedStoreDataQPreg_5 <= _T_2371[191:160];
    shiftedStoreDataQPreg_6 <= _T_2371[223:192];
    shiftedStoreDataQPreg_7 <= _T_2371[255:224];
    addrKnownPReg_0 <= addrKnown_0;
    addrKnownPReg_1 <= addrKnown_1;
    addrKnownPReg_2 <= addrKnown_2;
    addrKnownPReg_3 <= addrKnown_3;
    addrKnownPReg_4 <= addrKnown_4;
    addrKnownPReg_5 <= addrKnown_5;
    addrKnownPReg_6 <= addrKnown_6;
    addrKnownPReg_7 <= addrKnown_7;
    dataKnownPReg_0 <= dataKnown_0;
    dataKnownPReg_1 <= dataKnown_1;
    dataKnownPReg_2 <= dataKnown_2;
    dataKnownPReg_3 <= dataKnown_3;
    dataKnownPReg_4 <= dataKnown_4;
    dataKnownPReg_5 <= dataKnown_5;
    dataKnownPReg_6 <= dataKnown_6;
    dataKnownPReg_7 <= dataKnown_7;
    if (reset) begin
      prevPriorityRequest_7 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_7 <= priorityLoadRequest_7;
      end else begin
        prevPriorityRequest_7 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_6 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_6 <= priorityLoadRequest_6;
      end else begin
        prevPriorityRequest_6 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_5 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_5 <= priorityLoadRequest_5;
      end else begin
        prevPriorityRequest_5 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_4 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_4 <= priorityLoadRequest_4;
      end else begin
        prevPriorityRequest_4 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_3 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_3 <= priorityLoadRequest_3;
      end else begin
        prevPriorityRequest_3 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_2 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_2 <= priorityLoadRequest_2;
      end else begin
        prevPriorityRequest_2 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_1 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_1 <= priorityLoadRequest_1;
      end else begin
        prevPriorityRequest_1 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_0 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_0 <= priorityLoadRequest_0;
      end else begin
        prevPriorityRequest_0 <= 1'h0;
      end
    end
  end
endmodule
module GROUP_ALLOCATOR_LSQ_A( // @[:@12018.2]
  output [2:0] io_bbLoadOffsets_0, // @[:@12021.4]
  output [2:0] io_bbLoadOffsets_1, // @[:@12021.4]
  output [2:0] io_bbLoadOffsets_2, // @[:@12021.4]
  output [2:0] io_bbLoadOffsets_3, // @[:@12021.4]
  output [2:0] io_bbLoadOffsets_4, // @[:@12021.4]
  output [2:0] io_bbLoadOffsets_5, // @[:@12021.4]
  output [2:0] io_bbLoadOffsets_6, // @[:@12021.4]
  output [2:0] io_bbLoadOffsets_7, // @[:@12021.4]
  output       io_bbLoadPorts_1, // @[:@12021.4]
  output [1:0] io_bbNumLoads, // @[:@12021.4]
  input  [2:0] io_loadTail, // @[:@12021.4]
  input  [2:0] io_loadHead, // @[:@12021.4]
  input        io_loadEmpty, // @[:@12021.4]
  output [2:0] io_bbStoreOffsets_0, // @[:@12021.4]
  output [2:0] io_bbStoreOffsets_1, // @[:@12021.4]
  output [2:0] io_bbStoreOffsets_2, // @[:@12021.4]
  output [2:0] io_bbStoreOffsets_3, // @[:@12021.4]
  output [2:0] io_bbStoreOffsets_4, // @[:@12021.4]
  output [2:0] io_bbStoreOffsets_5, // @[:@12021.4]
  output [2:0] io_bbStoreOffsets_6, // @[:@12021.4]
  output [2:0] io_bbStoreOffsets_7, // @[:@12021.4]
  output       io_bbStorePorts_1, // @[:@12021.4]
  output [1:0] io_bbNumStores, // @[:@12021.4]
  input  [2:0] io_storeTail, // @[:@12021.4]
  input  [2:0] io_storeHead, // @[:@12021.4]
  input        io_storeEmpty, // @[:@12021.4]
  output       io_bbStart, // @[:@12021.4]
  input        io_bbStartSignals_0, // @[:@12021.4]
  output       io_readyToPrevious_0, // @[:@12021.4]
  output       io_loadPortsEnable_0, // @[:@12021.4]
  output       io_loadPortsEnable_1, // @[:@12021.4]
  output       io_storePortsEnable_0, // @[:@12021.4]
  output       io_storePortsEnable_1 // @[:@12021.4]
);
  wire  _T_180; // @[GroupAllocator.scala 42:25:@12024.4]
  wire  _T_181; // @[GroupAllocator.scala 42:16:@12025.4]
  wire [3:0] _GEN_36; // @[GroupAllocator.scala 43:36:@12027.6]
  wire [4:0] _T_183; // @[GroupAllocator.scala 43:36:@12027.6]
  wire [4:0] _T_184; // @[GroupAllocator.scala 43:36:@12028.6]
  wire [3:0] _T_185; // @[GroupAllocator.scala 43:36:@12029.6]
  wire [3:0] _GEN_37; // @[GroupAllocator.scala 43:43:@12030.6]
  wire [4:0] _T_186; // @[GroupAllocator.scala 43:43:@12030.6]
  wire [3:0] _T_187; // @[GroupAllocator.scala 43:43:@12031.6]
  wire [3:0] _T_188; // @[GroupAllocator.scala 45:22:@12035.6]
  wire [3:0] _T_189; // @[GroupAllocator.scala 45:22:@12036.6]
  wire [2:0] _T_190; // @[GroupAllocator.scala 45:22:@12037.6]
  wire [3:0] emptyLoadSlots; // @[GroupAllocator.scala 42:34:@12026.4]
  wire  _T_192; // @[GroupAllocator.scala 42:25:@12041.4]
  wire  _T_193; // @[GroupAllocator.scala 42:16:@12042.4]
  wire [3:0] _GEN_38; // @[GroupAllocator.scala 43:36:@12044.6]
  wire [4:0] _T_195; // @[GroupAllocator.scala 43:36:@12044.6]
  wire [4:0] _T_196; // @[GroupAllocator.scala 43:36:@12045.6]
  wire [3:0] _T_197; // @[GroupAllocator.scala 43:36:@12046.6]
  wire [3:0] _GEN_39; // @[GroupAllocator.scala 43:43:@12047.6]
  wire [4:0] _T_198; // @[GroupAllocator.scala 43:43:@12047.6]
  wire [3:0] _T_199; // @[GroupAllocator.scala 43:43:@12048.6]
  wire [3:0] _T_200; // @[GroupAllocator.scala 45:22:@12052.6]
  wire [3:0] _T_201; // @[GroupAllocator.scala 45:22:@12053.6]
  wire [2:0] _T_202; // @[GroupAllocator.scala 45:22:@12054.6]
  wire [3:0] emptyStoreSlots; // @[GroupAllocator.scala 42:34:@12043.4]
  wire  _T_204; // @[GroupAllocator.scala 54:19:@12057.4]
  wire  _T_206; // @[GroupAllocator.scala 54:50:@12058.4]
  wire [4:0] _T_493; // @[GroupAllocator.scala 110:34:@12222.6]
  wire [3:0] _T_494; // @[GroupAllocator.scala 110:34:@12223.6]
  wire [4:0] _T_496; // @[GroupAllocator.scala 110:55:@12224.6]
  wire [4:0] _T_497; // @[GroupAllocator.scala 110:55:@12225.6]
  wire [3:0] _T_498; // @[GroupAllocator.scala 110:55:@12226.6]
  wire [4:0] _T_500; // @[util.scala 10:8:@12227.6]
  wire [4:0] _GEN_0; // @[util.scala 10:14:@12228.6]
  wire [3:0] _T_501; // @[util.scala 10:14:@12228.6]
  wire [2:0] _T_504; // @[GroupAllocator.scala 110:90:@12229.6 GroupAllocator.scala 110:90:@12230.6]
  wire [4:0] _T_663; // @[GroupAllocator.scala 115:33:@12322.6]
  wire [3:0] _T_664; // @[GroupAllocator.scala 115:33:@12323.6]
  wire [4:0] _T_666; // @[GroupAllocator.scala 115:54:@12324.6]
  wire [4:0] _T_667; // @[GroupAllocator.scala 115:54:@12325.6]
  wire [3:0] _T_668; // @[GroupAllocator.scala 115:54:@12326.6]
  wire [4:0] _T_670; // @[util.scala 10:8:@12327.6]
  wire [4:0] _GEN_1; // @[util.scala 10:14:@12328.6]
  wire [3:0] _T_671; // @[util.scala 10:14:@12328.6]
  wire [4:0] _T_698; // @[util.scala 10:8:@12345.6]
  wire [4:0] _GEN_2; // @[util.scala 10:14:@12346.6]
  wire [3:0] _T_699; // @[util.scala 10:14:@12346.6]
  wire [2:0] _T_674; // @[GroupAllocator.scala 115:89:@12329.6 GroupAllocator.scala 115:89:@12330.6]
  wire [2:0] _T_702; // @[GroupAllocator.scala 115:89:@12347.6 GroupAllocator.scala 115:89:@12348.6]
  assign _T_180 = io_loadHead < io_loadTail; // @[GroupAllocator.scala 42:25:@12024.4]
  assign _T_181 = io_loadEmpty | _T_180; // @[GroupAllocator.scala 42:16:@12025.4]
  assign _GEN_36 = {{1'd0}, io_loadTail}; // @[GroupAllocator.scala 43:36:@12027.6]
  assign _T_183 = 4'h8 - _GEN_36; // @[GroupAllocator.scala 43:36:@12027.6]
  assign _T_184 = $unsigned(_T_183); // @[GroupAllocator.scala 43:36:@12028.6]
  assign _T_185 = _T_184[3:0]; // @[GroupAllocator.scala 43:36:@12029.6]
  assign _GEN_37 = {{1'd0}, io_loadHead}; // @[GroupAllocator.scala 43:43:@12030.6]
  assign _T_186 = _T_185 + _GEN_37; // @[GroupAllocator.scala 43:43:@12030.6]
  assign _T_187 = _T_185 + _GEN_37; // @[GroupAllocator.scala 43:43:@12031.6]
  assign _T_188 = io_loadHead - io_loadTail; // @[GroupAllocator.scala 45:22:@12035.6]
  assign _T_189 = $unsigned(_T_188); // @[GroupAllocator.scala 45:22:@12036.6]
  assign _T_190 = _T_189[2:0]; // @[GroupAllocator.scala 45:22:@12037.6]
  assign emptyLoadSlots = _T_181 ? _T_187 : {{1'd0}, _T_190}; // @[GroupAllocator.scala 42:34:@12026.4]
  assign _T_192 = io_storeHead < io_storeTail; // @[GroupAllocator.scala 42:25:@12041.4]
  assign _T_193 = io_storeEmpty | _T_192; // @[GroupAllocator.scala 42:16:@12042.4]
  assign _GEN_38 = {{1'd0}, io_storeTail}; // @[GroupAllocator.scala 43:36:@12044.6]
  assign _T_195 = 4'h8 - _GEN_38; // @[GroupAllocator.scala 43:36:@12044.6]
  assign _T_196 = $unsigned(_T_195); // @[GroupAllocator.scala 43:36:@12045.6]
  assign _T_197 = _T_196[3:0]; // @[GroupAllocator.scala 43:36:@12046.6]
  assign _GEN_39 = {{1'd0}, io_storeHead}; // @[GroupAllocator.scala 43:43:@12047.6]
  assign _T_198 = _T_197 + _GEN_39; // @[GroupAllocator.scala 43:43:@12047.6]
  assign _T_199 = _T_197 + _GEN_39; // @[GroupAllocator.scala 43:43:@12048.6]
  assign _T_200 = io_storeHead - io_storeTail; // @[GroupAllocator.scala 45:22:@12052.6]
  assign _T_201 = $unsigned(_T_200); // @[GroupAllocator.scala 45:22:@12053.6]
  assign _T_202 = _T_201[2:0]; // @[GroupAllocator.scala 45:22:@12054.6]
  assign emptyStoreSlots = _T_193 ? _T_199 : {{1'd0}, _T_202}; // @[GroupAllocator.scala 42:34:@12043.4]
  assign _T_204 = 4'h2 <= emptyStoreSlots; // @[GroupAllocator.scala 54:19:@12057.4]
  assign _T_206 = 4'h2 <= emptyLoadSlots; // @[GroupAllocator.scala 54:50:@12058.4]
  assign _T_493 = _GEN_38 + 4'h8; // @[GroupAllocator.scala 110:34:@12222.6]
  assign _T_494 = _GEN_38 + 4'h8; // @[GroupAllocator.scala 110:34:@12223.6]
  assign _T_496 = _T_494 - 4'h1; // @[GroupAllocator.scala 110:55:@12224.6]
  assign _T_497 = $unsigned(_T_496); // @[GroupAllocator.scala 110:55:@12225.6]
  assign _T_498 = _T_497[3:0]; // @[GroupAllocator.scala 110:55:@12226.6]
  assign _T_500 = {{1'd0}, _T_498}; // @[util.scala 10:8:@12227.6]
  assign _GEN_0 = _T_500 % 5'h8; // @[util.scala 10:14:@12228.6]
  assign _T_501 = _GEN_0[3:0]; // @[util.scala 10:14:@12228.6]
  assign _T_504 = _T_501[2:0]; // @[GroupAllocator.scala 110:90:@12229.6 GroupAllocator.scala 110:90:@12230.6]
  assign _T_663 = _GEN_36 + 4'h8; // @[GroupAllocator.scala 115:33:@12322.6]
  assign _T_664 = _GEN_36 + 4'h8; // @[GroupAllocator.scala 115:33:@12323.6]
  assign _T_666 = _T_664 - 4'h1; // @[GroupAllocator.scala 115:54:@12324.6]
  assign _T_667 = $unsigned(_T_666); // @[GroupAllocator.scala 115:54:@12325.6]
  assign _T_668 = _T_667[3:0]; // @[GroupAllocator.scala 115:54:@12326.6]
  assign _T_670 = 4'h2 + _T_668; // @[util.scala 10:8:@12327.6]
  assign _GEN_1 = _T_670 % 5'h8; // @[util.scala 10:14:@12328.6]
  assign _T_671 = _GEN_1[3:0]; // @[util.scala 10:14:@12328.6]
  assign _T_698 = {{1'd0}, _T_668}; // @[util.scala 10:8:@12345.6]
  assign _GEN_2 = _T_698 % 5'h8; // @[util.scala 10:14:@12346.6]
  assign _T_699 = _GEN_2[3:0]; // @[util.scala 10:14:@12346.6]
  assign _T_674 = _T_671[2:0]; // @[GroupAllocator.scala 115:89:@12329.6 GroupAllocator.scala 115:89:@12330.6]
  assign _T_702 = _T_699[2:0]; // @[GroupAllocator.scala 115:89:@12347.6 GroupAllocator.scala 115:89:@12348.6]
  assign io_bbLoadOffsets_0 = io_bbStart ? _T_504 : 3'h0; // @[GroupAllocator.scala 89:20:@12125.4 GroupAllocator.scala 106:22:@12305.6]
  assign io_bbLoadOffsets_1 = io_bbStart ? _T_504 : 3'h0; // @[GroupAllocator.scala 89:20:@12126.4 GroupAllocator.scala 106:22:@12306.6]
  assign io_bbLoadOffsets_2 = io_bbStart ? _T_504 : 3'h0; // @[GroupAllocator.scala 89:20:@12127.4 GroupAllocator.scala 106:22:@12307.6]
  assign io_bbLoadOffsets_3 = io_bbStart ? _T_504 : 3'h0; // @[GroupAllocator.scala 89:20:@12128.4 GroupAllocator.scala 106:22:@12308.6]
  assign io_bbLoadOffsets_4 = io_bbStart ? _T_504 : 3'h0; // @[GroupAllocator.scala 89:20:@12129.4 GroupAllocator.scala 106:22:@12309.6]
  assign io_bbLoadOffsets_5 = io_bbStart ? _T_504 : 3'h0; // @[GroupAllocator.scala 89:20:@12130.4 GroupAllocator.scala 106:22:@12310.6]
  assign io_bbLoadOffsets_6 = io_bbStart ? _T_504 : 3'h0; // @[GroupAllocator.scala 89:20:@12131.4 GroupAllocator.scala 106:22:@12311.6]
  assign io_bbLoadOffsets_7 = io_bbStart ? _T_504 : 3'h0; // @[GroupAllocator.scala 89:20:@12132.4 GroupAllocator.scala 106:22:@12312.6]
  assign io_bbLoadPorts_1 = io_bbStart; // @[GroupAllocator.scala 87:18:@12092.4 GroupAllocator.scala 95:20:@12178.6]
  assign io_bbNumLoads = io_bbStart ? 2'h2 : 2'h0; // @[GroupAllocator.scala 85:17:@12080.4 GroupAllocator.scala 93:19:@12153.6]
  assign io_bbStoreOffsets_0 = io_bbStart ? _T_674 : 3'h0; // @[GroupAllocator.scala 90:21:@12142.4 GroupAllocator.scala 111:23:@12405.6]
  assign io_bbStoreOffsets_1 = io_bbStart ? _T_674 : 3'h0; // @[GroupAllocator.scala 90:21:@12143.4 GroupAllocator.scala 111:23:@12406.6]
  assign io_bbStoreOffsets_2 = io_bbStart ? _T_702 : 3'h0; // @[GroupAllocator.scala 90:21:@12144.4 GroupAllocator.scala 111:23:@12407.6]
  assign io_bbStoreOffsets_3 = io_bbStart ? _T_702 : 3'h0; // @[GroupAllocator.scala 90:21:@12145.4 GroupAllocator.scala 111:23:@12408.6]
  assign io_bbStoreOffsets_4 = io_bbStart ? _T_702 : 3'h0; // @[GroupAllocator.scala 90:21:@12146.4 GroupAllocator.scala 111:23:@12409.6]
  assign io_bbStoreOffsets_5 = io_bbStart ? _T_702 : 3'h0; // @[GroupAllocator.scala 90:21:@12147.4 GroupAllocator.scala 111:23:@12410.6]
  assign io_bbStoreOffsets_6 = io_bbStart ? _T_702 : 3'h0; // @[GroupAllocator.scala 90:21:@12148.4 GroupAllocator.scala 111:23:@12411.6]
  assign io_bbStoreOffsets_7 = io_bbStart ? _T_702 : 3'h0; // @[GroupAllocator.scala 90:21:@12149.4 GroupAllocator.scala 111:23:@12412.6]
  assign io_bbStorePorts_1 = io_bbStart; // @[GroupAllocator.scala 88:19:@12109.4 GroupAllocator.scala 100:21:@12206.6]
  assign io_bbNumStores = io_bbStart ? 2'h2 : 2'h0; // @[GroupAllocator.scala 86:18:@12081.4 GroupAllocator.scala 94:20:@12156.6]
  assign io_bbStart = io_readyToPrevious_0 & io_bbStartSignals_0; // @[GroupAllocator.scala 59:14:@12067.4]
  assign io_readyToPrevious_0 = _T_204 & _T_206; // @[GroupAllocator.scala 53:22:@12062.4]
  assign io_loadPortsEnable_0 = io_bbStart; // @[GroupAllocator.scala 69:29:@12070.4]
  assign io_loadPortsEnable_1 = io_bbStart; // @[GroupAllocator.scala 69:29:@12073.4]
  assign io_storePortsEnable_0 = io_bbStart; // @[GroupAllocator.scala 78:30:@12076.4]
  assign io_storePortsEnable_1 = io_bbStart; // @[GroupAllocator.scala 78:30:@12079.4]
endmodule
module LOAD_PORT_LSQ_A( // @[:@12415.2]
  input         clock, // @[:@12416.4]
  input         reset, // @[:@12417.4]
  output        io_addrFromPrev_ready, // @[:@12418.4]
  input         io_addrFromPrev_valid, // @[:@12418.4]
  input  [31:0] io_addrFromPrev_bits, // @[:@12418.4]
  input         io_portEnable, // @[:@12418.4]
  input         io_dataToNext_ready, // @[:@12418.4]
  output        io_dataToNext_valid, // @[:@12418.4]
  output [31:0] io_dataToNext_bits, // @[:@12418.4]
  output        io_loadAddrEnable, // @[:@12418.4]
  output [31:0] io_addrToLoadQueue, // @[:@12418.4]
  output        io_dataFromLoadQueue_ready, // @[:@12418.4]
  input         io_dataFromLoadQueue_valid, // @[:@12418.4]
  input  [31:0] io_dataFromLoadQueue_bits // @[:@12418.4]
);
  reg [3:0] cnt; // @[LoadPort.scala 23:20:@12420.4]
  reg [31:0] _RAND_0;
  wire  _T_44; // @[LoadPort.scala 26:25:@12421.4]
  wire  _T_45; // @[LoadPort.scala 26:22:@12422.4]
  wire  _T_47; // @[LoadPort.scala 26:51:@12423.4]
  wire  _T_48; // @[LoadPort.scala 26:44:@12424.4]
  wire [4:0] _T_50; // @[LoadPort.scala 27:16:@12426.6]
  wire [3:0] _T_51; // @[LoadPort.scala 27:16:@12427.6]
  wire  _T_53; // @[LoadPort.scala 28:35:@12431.6]
  wire  _T_54; // @[LoadPort.scala 28:32:@12432.6]
  wire  _T_56; // @[LoadPort.scala 28:57:@12433.6]
  wire  _T_57; // @[LoadPort.scala 28:50:@12434.6]
  wire [4:0] _T_59; // @[LoadPort.scala 29:16:@12436.8]
  wire [4:0] _T_60; // @[LoadPort.scala 29:16:@12437.8]
  wire [3:0] _T_61; // @[LoadPort.scala 29:16:@12438.8]
  wire [3:0] _GEN_0; // @[LoadPort.scala 28:66:@12435.6]
  wire [3:0] _GEN_1; // @[LoadPort.scala 26:75:@12425.4]
  wire  _T_63; // @[LoadPort.scala 33:28:@12442.4]
  assign _T_44 = io_loadAddrEnable == 1'h0; // @[LoadPort.scala 26:25:@12421.4]
  assign _T_45 = io_portEnable & _T_44; // @[LoadPort.scala 26:22:@12422.4]
  assign _T_47 = cnt != 4'h8; // @[LoadPort.scala 26:51:@12423.4]
  assign _T_48 = _T_45 & _T_47; // @[LoadPort.scala 26:44:@12424.4]
  assign _T_50 = cnt + 4'h1; // @[LoadPort.scala 27:16:@12426.6]
  assign _T_51 = cnt + 4'h1; // @[LoadPort.scala 27:16:@12427.6]
  assign _T_53 = io_portEnable == 1'h0; // @[LoadPort.scala 28:35:@12431.6]
  assign _T_54 = io_loadAddrEnable & _T_53; // @[LoadPort.scala 28:32:@12432.6]
  assign _T_56 = cnt != 4'h0; // @[LoadPort.scala 28:57:@12433.6]
  assign _T_57 = _T_54 & _T_56; // @[LoadPort.scala 28:50:@12434.6]
  assign _T_59 = cnt - 4'h1; // @[LoadPort.scala 29:16:@12436.8]
  assign _T_60 = $unsigned(_T_59); // @[LoadPort.scala 29:16:@12437.8]
  assign _T_61 = _T_60[3:0]; // @[LoadPort.scala 29:16:@12438.8]
  assign _GEN_0 = _T_57 ? _T_61 : cnt; // @[LoadPort.scala 28:66:@12435.6]
  assign _GEN_1 = _T_48 ? _T_51 : _GEN_0; // @[LoadPort.scala 26:75:@12425.4]
  assign _T_63 = cnt > 4'h0; // @[LoadPort.scala 33:28:@12442.4]
  assign io_addrFromPrev_ready = cnt > 4'h0; // @[LoadPort.scala 34:25:@12446.4]
  assign io_dataToNext_valid = io_dataFromLoadQueue_valid; // @[LoadPort.scala 35:17:@12448.4]
  assign io_dataToNext_bits = io_dataFromLoadQueue_bits; // @[LoadPort.scala 35:17:@12447.4]
  assign io_loadAddrEnable = _T_63 & io_addrFromPrev_valid; // @[LoadPort.scala 33:21:@12444.4]
  assign io_addrToLoadQueue = io_addrFromPrev_bits; // @[LoadPort.scala 32:22:@12441.4]
  assign io_dataFromLoadQueue_ready = io_dataToNext_ready; // @[LoadPort.scala 35:17:@12449.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 4'h0;
    end else begin
      if (_T_48) begin
        cnt <= _T_51;
      end else begin
        if (_T_57) begin
          cnt <= _T_61;
        end
      end
    end
  end
endmodule
module STORE_DATA_PORT_LSQ_A( // @[:@12487.2]
  input         clock, // @[:@12488.4]
  input         reset, // @[:@12489.4]
  output        io_dataFromPrev_ready, // @[:@12490.4]
  input         io_dataFromPrev_valid, // @[:@12490.4]
  input  [31:0] io_dataFromPrev_bits, // @[:@12490.4]
  input         io_portEnable, // @[:@12490.4]
  output        io_storeDataEnable, // @[:@12490.4]
  output [31:0] io_dataToStoreQueue // @[:@12490.4]
);
  reg [3:0] cnt; // @[StoreDataPort.scala 21:20:@12492.4]
  reg [31:0] _RAND_0;
  wire  _T_26; // @[StoreDataPort.scala 24:25:@12493.4]
  wire  _T_27; // @[StoreDataPort.scala 24:22:@12494.4]
  wire  _T_29; // @[StoreDataPort.scala 24:52:@12495.4]
  wire  _T_30; // @[StoreDataPort.scala 24:45:@12496.4]
  wire [4:0] _T_32; // @[StoreDataPort.scala 25:16:@12498.6]
  wire [3:0] _T_33; // @[StoreDataPort.scala 25:16:@12499.6]
  wire  _T_35; // @[StoreDataPort.scala 26:36:@12503.6]
  wire  _T_36; // @[StoreDataPort.scala 26:33:@12504.6]
  wire  _T_38; // @[StoreDataPort.scala 26:58:@12505.6]
  wire  _T_39; // @[StoreDataPort.scala 26:51:@12506.6]
  wire [4:0] _T_41; // @[StoreDataPort.scala 27:16:@12508.8]
  wire [4:0] _T_42; // @[StoreDataPort.scala 27:16:@12509.8]
  wire [3:0] _T_43; // @[StoreDataPort.scala 27:16:@12510.8]
  wire [3:0] _GEN_0; // @[StoreDataPort.scala 26:67:@12507.6]
  wire [3:0] _GEN_1; // @[StoreDataPort.scala 24:76:@12497.4]
  wire  _T_45; // @[StoreDataPort.scala 31:29:@12514.4]
  assign _T_26 = io_storeDataEnable == 1'h0; // @[StoreDataPort.scala 24:25:@12493.4]
  assign _T_27 = io_portEnable & _T_26; // @[StoreDataPort.scala 24:22:@12494.4]
  assign _T_29 = cnt != 4'h8; // @[StoreDataPort.scala 24:52:@12495.4]
  assign _T_30 = _T_27 & _T_29; // @[StoreDataPort.scala 24:45:@12496.4]
  assign _T_32 = cnt + 4'h1; // @[StoreDataPort.scala 25:16:@12498.6]
  assign _T_33 = cnt + 4'h1; // @[StoreDataPort.scala 25:16:@12499.6]
  assign _T_35 = io_portEnable == 1'h0; // @[StoreDataPort.scala 26:36:@12503.6]
  assign _T_36 = io_storeDataEnable & _T_35; // @[StoreDataPort.scala 26:33:@12504.6]
  assign _T_38 = cnt != 4'h0; // @[StoreDataPort.scala 26:58:@12505.6]
  assign _T_39 = _T_36 & _T_38; // @[StoreDataPort.scala 26:51:@12506.6]
  assign _T_41 = cnt - 4'h1; // @[StoreDataPort.scala 27:16:@12508.8]
  assign _T_42 = $unsigned(_T_41); // @[StoreDataPort.scala 27:16:@12509.8]
  assign _T_43 = _T_42[3:0]; // @[StoreDataPort.scala 27:16:@12510.8]
  assign _GEN_0 = _T_39 ? _T_43 : cnt; // @[StoreDataPort.scala 26:67:@12507.6]
  assign _GEN_1 = _T_30 ? _T_33 : _GEN_0; // @[StoreDataPort.scala 24:76:@12497.4]
  assign _T_45 = cnt > 4'h0; // @[StoreDataPort.scala 31:29:@12514.4]
  assign io_dataFromPrev_ready = cnt > 4'h0; // @[StoreDataPort.scala 32:25:@12518.4]
  assign io_storeDataEnable = _T_45 & io_dataFromPrev_valid; // @[StoreDataPort.scala 31:22:@12516.4]
  assign io_dataToStoreQueue = io_dataFromPrev_bits; // @[StoreDataPort.scala 30:23:@12513.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 4'h0;
    end else begin
      if (_T_30) begin
        cnt <= _T_33;
      end else begin
        if (_T_39) begin
          cnt <= _T_43;
        end
      end
    end
  end
endmodule
module LSQ_A( // @[:@12619.2]
  input         clock, // @[:@12620.4]
  input         reset, // @[:@12621.4]
  output [31:0] io_storeDataOut, // @[:@12622.4]
  output [31:0] io_storeAddrOut, // @[:@12622.4]
  output        io_storeEnable, // @[:@12622.4]
  input         io_memIsReadyForStores, // @[:@12622.4]
  input  [31:0] io_loadDataIn, // @[:@12622.4]
  output [31:0] io_loadAddrOut, // @[:@12622.4]
  output        io_loadEnable, // @[:@12622.4]
  input         io_memIsReadyForLoads, // @[:@12622.4]
  input         io_bbpValids_0, // @[:@12622.4]
  output        io_bbReadyToPrevs_0, // @[:@12622.4]
  output        io_rdPortsPrev_0_ready, // @[:@12622.4]
  input         io_rdPortsPrev_0_valid, // @[:@12622.4]
  input  [31:0] io_rdPortsPrev_0_bits, // @[:@12622.4]
  output        io_rdPortsPrev_1_ready, // @[:@12622.4]
  input         io_rdPortsPrev_1_valid, // @[:@12622.4]
  input  [31:0] io_rdPortsPrev_1_bits, // @[:@12622.4]
  input         io_rdPortsNext_0_ready, // @[:@12622.4]
  output        io_rdPortsNext_0_valid, // @[:@12622.4]
  output [31:0] io_rdPortsNext_0_bits, // @[:@12622.4]
  input         io_rdPortsNext_1_ready, // @[:@12622.4]
  output        io_rdPortsNext_1_valid, // @[:@12622.4]
  output [31:0] io_rdPortsNext_1_bits, // @[:@12622.4]
  output        io_wrAddrPorts_0_ready, // @[:@12622.4]
  input         io_wrAddrPorts_0_valid, // @[:@12622.4]
  input  [31:0] io_wrAddrPorts_0_bits, // @[:@12622.4]
  output        io_wrAddrPorts_1_ready, // @[:@12622.4]
  input         io_wrAddrPorts_1_valid, // @[:@12622.4]
  input  [31:0] io_wrAddrPorts_1_bits, // @[:@12622.4]
  output        io_wrDataPorts_0_ready, // @[:@12622.4]
  input         io_wrDataPorts_0_valid, // @[:@12622.4]
  input  [31:0] io_wrDataPorts_0_bits, // @[:@12622.4]
  output        io_wrDataPorts_1_ready, // @[:@12622.4]
  input         io_wrDataPorts_1_valid, // @[:@12622.4]
  input  [31:0] io_wrDataPorts_1_bits, // @[:@12622.4]
  output        io_Empty_Valid // @[:@12622.4]
);
  wire  storeQ_clock; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_reset; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_bbStart; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_bbStoreOffsets_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_bbStoreOffsets_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_bbStoreOffsets_2; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_bbStoreOffsets_3; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_bbStoreOffsets_4; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_bbStoreOffsets_5; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_bbStoreOffsets_6; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_bbStoreOffsets_7; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_bbStorePorts_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [1:0] storeQ_io_bbNumStores; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_storeTail; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_storeHead; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeEmpty; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_loadTail; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [2:0] storeQ_io_loadHead; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadEmpty; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadAddressDone_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadAddressDone_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadAddressDone_2; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadAddressDone_3; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadAddressDone_4; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadAddressDone_5; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadAddressDone_6; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadAddressDone_7; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadDataDone_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadDataDone_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadDataDone_2; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadDataDone_3; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadDataDone_4; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadDataDone_5; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadDataDone_6; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_loadDataDone_7; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_loadAddressQueue_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_loadAddressQueue_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_loadAddressQueue_2; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_loadAddressQueue_3; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_loadAddressQueue_4; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_loadAddressQueue_5; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_loadAddressQueue_6; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_loadAddressQueue_7; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataEnable_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeDataEnable_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_dataFromStorePorts_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_dataFromStorePorts_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrEnable_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeAddrEnable_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_addressFromStorePorts_0; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_addressFromStorePorts_1; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 72:22:@12653.4]
  wire [31:0] storeQ_io_storeDataToMem; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  storeQ_io_memIsReadyForStores; // @[LSQBRAM.scala 72:22:@12653.4]
  wire  loadQ_clock; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_reset; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_bbStart; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_bbLoadOffsets_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_bbLoadOffsets_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_bbLoadOffsets_2; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_bbLoadOffsets_3; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_bbLoadOffsets_4; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_bbLoadOffsets_5; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_bbLoadOffsets_6; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_bbLoadOffsets_7; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_bbLoadPorts_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [1:0] loadQ_io_bbNumLoads; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_loadTail; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_loadHead; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadEmpty; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_storeTail; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] loadQ_io_storeHead; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeEmpty; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeAddrDone_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeAddrDone_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeAddrDone_2; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeAddrDone_3; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeAddrDone_4; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeAddrDone_5; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeAddrDone_6; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeAddrDone_7; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeDataDone_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeDataDone_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeDataDone_2; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeDataDone_3; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeDataDone_4; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeDataDone_5; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeDataDone_6; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_storeDataDone_7; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeDataQueue_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeDataQueue_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeDataQueue_2; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeDataQueue_3; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeDataQueue_4; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeDataQueue_5; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeDataQueue_6; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_storeDataQueue_7; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrEnable_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadAddrEnable_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_0; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_1; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadPorts_0_ready; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadPorts_1_ready; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadPorts_1_valid; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadPorts_1_bits; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadDataFromMem; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [31:0] loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 73:21:@12656.4]
  wire  loadQ_io_memIsReadyForLoads; // @[LSQBRAM.scala 73:21:@12656.4]
  wire [2:0] GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_bbLoadPorts_1; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [1:0] GA_io_bbNumLoads; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_loadTail; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_loadHead; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_loadEmpty; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_bbStorePorts_1; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [1:0] GA_io_bbNumStores; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_storeTail; // @[LSQBRAM.scala 74:18:@12659.4]
  wire [2:0] GA_io_storeHead; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_storeEmpty; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_bbStart; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_bbStartSignals_0; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_readyToPrevious_0; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_loadPortsEnable_1; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_storePortsEnable_0; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  GA_io_storePortsEnable_1; // @[LSQBRAM.scala 74:18:@12659.4]
  wire  LOAD_PORT_LSQ_A_clock; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_reset; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@12662.4]
  wire [31:0] LOAD_PORT_LSQ_A_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_io_portEnable; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@12662.4]
  wire [31:0] LOAD_PORT_LSQ_A_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@12662.4]
  wire [31:0] LOAD_PORT_LSQ_A_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@12662.4]
  wire [31:0] LOAD_PORT_LSQ_A_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@12662.4]
  wire  LOAD_PORT_LSQ_A_1_clock; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  LOAD_PORT_LSQ_A_1_reset; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  LOAD_PORT_LSQ_A_1_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  LOAD_PORT_LSQ_A_1_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@12665.4]
  wire [31:0] LOAD_PORT_LSQ_A_1_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  LOAD_PORT_LSQ_A_1_io_portEnable; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  LOAD_PORT_LSQ_A_1_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  LOAD_PORT_LSQ_A_1_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@12665.4]
  wire [31:0] LOAD_PORT_LSQ_A_1_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  LOAD_PORT_LSQ_A_1_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@12665.4]
  wire [31:0] LOAD_PORT_LSQ_A_1_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  LOAD_PORT_LSQ_A_1_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  LOAD_PORT_LSQ_A_1_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@12665.4]
  wire [31:0] LOAD_PORT_LSQ_A_1_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@12665.4]
  wire  STORE_DATA_PORT_LSQ_A_clock; // @[LSQBRAM.scala 80:11:@12693.4]
  wire  STORE_DATA_PORT_LSQ_A_reset; // @[LSQBRAM.scala 80:11:@12693.4]
  wire  STORE_DATA_PORT_LSQ_A_io_dataFromPrev_ready; // @[LSQBRAM.scala 80:11:@12693.4]
  wire  STORE_DATA_PORT_LSQ_A_io_dataFromPrev_valid; // @[LSQBRAM.scala 80:11:@12693.4]
  wire [31:0] STORE_DATA_PORT_LSQ_A_io_dataFromPrev_bits; // @[LSQBRAM.scala 80:11:@12693.4]
  wire  STORE_DATA_PORT_LSQ_A_io_portEnable; // @[LSQBRAM.scala 80:11:@12693.4]
  wire  STORE_DATA_PORT_LSQ_A_io_storeDataEnable; // @[LSQBRAM.scala 80:11:@12693.4]
  wire [31:0] STORE_DATA_PORT_LSQ_A_io_dataToStoreQueue; // @[LSQBRAM.scala 80:11:@12693.4]
  wire  STORE_DATA_PORT_LSQ_A_1_clock; // @[LSQBRAM.scala 80:11:@12696.4]
  wire  STORE_DATA_PORT_LSQ_A_1_reset; // @[LSQBRAM.scala 80:11:@12696.4]
  wire  STORE_DATA_PORT_LSQ_A_1_io_dataFromPrev_ready; // @[LSQBRAM.scala 80:11:@12696.4]
  wire  STORE_DATA_PORT_LSQ_A_1_io_dataFromPrev_valid; // @[LSQBRAM.scala 80:11:@12696.4]
  wire [31:0] STORE_DATA_PORT_LSQ_A_1_io_dataFromPrev_bits; // @[LSQBRAM.scala 80:11:@12696.4]
  wire  STORE_DATA_PORT_LSQ_A_1_io_portEnable; // @[LSQBRAM.scala 80:11:@12696.4]
  wire  STORE_DATA_PORT_LSQ_A_1_io_storeDataEnable; // @[LSQBRAM.scala 80:11:@12696.4]
  wire [31:0] STORE_DATA_PORT_LSQ_A_1_io_dataToStoreQueue; // @[LSQBRAM.scala 80:11:@12696.4]
  wire  STORE_ADDR_PORT_LSQ_A_clock; // @[LSQBRAM.scala 83:11:@12712.4]
  wire  STORE_ADDR_PORT_LSQ_A_reset; // @[LSQBRAM.scala 83:11:@12712.4]
  wire  STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_ready; // @[LSQBRAM.scala 83:11:@12712.4]
  wire  STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_valid; // @[LSQBRAM.scala 83:11:@12712.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_bits; // @[LSQBRAM.scala 83:11:@12712.4]
  wire  STORE_ADDR_PORT_LSQ_A_io_portEnable; // @[LSQBRAM.scala 83:11:@12712.4]
  wire  STORE_ADDR_PORT_LSQ_A_io_storeDataEnable; // @[LSQBRAM.scala 83:11:@12712.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_A_io_dataToStoreQueue; // @[LSQBRAM.scala 83:11:@12712.4]
  wire  STORE_ADDR_PORT_LSQ_A_1_clock; // @[LSQBRAM.scala 83:11:@12715.4]
  wire  STORE_ADDR_PORT_LSQ_A_1_reset; // @[LSQBRAM.scala 83:11:@12715.4]
  wire  STORE_ADDR_PORT_LSQ_A_1_io_dataFromPrev_ready; // @[LSQBRAM.scala 83:11:@12715.4]
  wire  STORE_ADDR_PORT_LSQ_A_1_io_dataFromPrev_valid; // @[LSQBRAM.scala 83:11:@12715.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_A_1_io_dataFromPrev_bits; // @[LSQBRAM.scala 83:11:@12715.4]
  wire  STORE_ADDR_PORT_LSQ_A_1_io_portEnable; // @[LSQBRAM.scala 83:11:@12715.4]
  wire  STORE_ADDR_PORT_LSQ_A_1_io_storeDataEnable; // @[LSQBRAM.scala 83:11:@12715.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_A_1_io_dataToStoreQueue; // @[LSQBRAM.scala 83:11:@12715.4]
  wire  storeEmpty; // @[LSQBRAM.scala 46:24:@12629.4 LSQBRAM.scala 151:14:@12921.4]
  wire  loadEmpty; // @[LSQBRAM.scala 52:23:@12635.4 LSQBRAM.scala 119:13:@12835.4]
  wire [7:0] storeTail; // @[LSQBRAM.scala 44:23:@12627.4 LSQBRAM.scala 149:13:@12919.4]
  wire [7:0] storeHead; // @[LSQBRAM.scala 45:23:@12628.4 LSQBRAM.scala 150:13:@12920.4]
  wire [7:0] loadTail; // @[LSQBRAM.scala 50:22:@12633.4 LSQBRAM.scala 117:12:@12833.4]
  wire [7:0] loadHead; // @[LSQBRAM.scala 51:22:@12634.4 LSQBRAM.scala 118:12:@12834.4]
  STORE_QUEUE_LSQ_A storeQ ( // @[LSQBRAM.scala 72:22:@12653.4]
    .clock(storeQ_clock),
    .reset(storeQ_reset),
    .io_bbStart(storeQ_io_bbStart),
    .io_bbStoreOffsets_0(storeQ_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(storeQ_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(storeQ_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(storeQ_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(storeQ_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(storeQ_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(storeQ_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(storeQ_io_bbStoreOffsets_7),
    .io_bbStorePorts_1(storeQ_io_bbStorePorts_1),
    .io_bbNumStores(storeQ_io_bbNumStores),
    .io_storeTail(storeQ_io_storeTail),
    .io_storeHead(storeQ_io_storeHead),
    .io_storeEmpty(storeQ_io_storeEmpty),
    .io_loadTail(storeQ_io_loadTail),
    .io_loadHead(storeQ_io_loadHead),
    .io_loadEmpty(storeQ_io_loadEmpty),
    .io_loadAddressDone_0(storeQ_io_loadAddressDone_0),
    .io_loadAddressDone_1(storeQ_io_loadAddressDone_1),
    .io_loadAddressDone_2(storeQ_io_loadAddressDone_2),
    .io_loadAddressDone_3(storeQ_io_loadAddressDone_3),
    .io_loadAddressDone_4(storeQ_io_loadAddressDone_4),
    .io_loadAddressDone_5(storeQ_io_loadAddressDone_5),
    .io_loadAddressDone_6(storeQ_io_loadAddressDone_6),
    .io_loadAddressDone_7(storeQ_io_loadAddressDone_7),
    .io_loadDataDone_0(storeQ_io_loadDataDone_0),
    .io_loadDataDone_1(storeQ_io_loadDataDone_1),
    .io_loadDataDone_2(storeQ_io_loadDataDone_2),
    .io_loadDataDone_3(storeQ_io_loadDataDone_3),
    .io_loadDataDone_4(storeQ_io_loadDataDone_4),
    .io_loadDataDone_5(storeQ_io_loadDataDone_5),
    .io_loadDataDone_6(storeQ_io_loadDataDone_6),
    .io_loadDataDone_7(storeQ_io_loadDataDone_7),
    .io_loadAddressQueue_0(storeQ_io_loadAddressQueue_0),
    .io_loadAddressQueue_1(storeQ_io_loadAddressQueue_1),
    .io_loadAddressQueue_2(storeQ_io_loadAddressQueue_2),
    .io_loadAddressQueue_3(storeQ_io_loadAddressQueue_3),
    .io_loadAddressQueue_4(storeQ_io_loadAddressQueue_4),
    .io_loadAddressQueue_5(storeQ_io_loadAddressQueue_5),
    .io_loadAddressQueue_6(storeQ_io_loadAddressQueue_6),
    .io_loadAddressQueue_7(storeQ_io_loadAddressQueue_7),
    .io_storeAddrDone_0(storeQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(storeQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(storeQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(storeQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(storeQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(storeQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(storeQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(storeQ_io_storeAddrDone_7),
    .io_storeDataDone_0(storeQ_io_storeDataDone_0),
    .io_storeDataDone_1(storeQ_io_storeDataDone_1),
    .io_storeDataDone_2(storeQ_io_storeDataDone_2),
    .io_storeDataDone_3(storeQ_io_storeDataDone_3),
    .io_storeDataDone_4(storeQ_io_storeDataDone_4),
    .io_storeDataDone_5(storeQ_io_storeDataDone_5),
    .io_storeDataDone_6(storeQ_io_storeDataDone_6),
    .io_storeDataDone_7(storeQ_io_storeDataDone_7),
    .io_storeAddrQueue_0(storeQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(storeQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(storeQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(storeQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(storeQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(storeQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(storeQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(storeQ_io_storeAddrQueue_7),
    .io_storeDataQueue_0(storeQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(storeQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(storeQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(storeQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(storeQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(storeQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(storeQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(storeQ_io_storeDataQueue_7),
    .io_storeDataEnable_0(storeQ_io_storeDataEnable_0),
    .io_storeDataEnable_1(storeQ_io_storeDataEnable_1),
    .io_dataFromStorePorts_0(storeQ_io_dataFromStorePorts_0),
    .io_dataFromStorePorts_1(storeQ_io_dataFromStorePorts_1),
    .io_storeAddrEnable_0(storeQ_io_storeAddrEnable_0),
    .io_storeAddrEnable_1(storeQ_io_storeAddrEnable_1),
    .io_addressFromStorePorts_0(storeQ_io_addressFromStorePorts_0),
    .io_addressFromStorePorts_1(storeQ_io_addressFromStorePorts_1),
    .io_storeAddrToMem(storeQ_io_storeAddrToMem),
    .io_storeDataToMem(storeQ_io_storeDataToMem),
    .io_storeEnableToMem(storeQ_io_storeEnableToMem),
    .io_memIsReadyForStores(storeQ_io_memIsReadyForStores)
  );
  LOAD_QUEUE_LSQ_A loadQ ( // @[LSQBRAM.scala 73:21:@12656.4]
    .clock(loadQ_clock),
    .reset(loadQ_reset),
    .io_bbStart(loadQ_io_bbStart),
    .io_bbLoadOffsets_0(loadQ_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(loadQ_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(loadQ_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(loadQ_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(loadQ_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(loadQ_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(loadQ_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(loadQ_io_bbLoadOffsets_7),
    .io_bbLoadPorts_1(loadQ_io_bbLoadPorts_1),
    .io_bbNumLoads(loadQ_io_bbNumLoads),
    .io_loadTail(loadQ_io_loadTail),
    .io_loadHead(loadQ_io_loadHead),
    .io_loadEmpty(loadQ_io_loadEmpty),
    .io_storeTail(loadQ_io_storeTail),
    .io_storeHead(loadQ_io_storeHead),
    .io_storeEmpty(loadQ_io_storeEmpty),
    .io_storeAddrDone_0(loadQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(loadQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(loadQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(loadQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(loadQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(loadQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(loadQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(loadQ_io_storeAddrDone_7),
    .io_storeDataDone_0(loadQ_io_storeDataDone_0),
    .io_storeDataDone_1(loadQ_io_storeDataDone_1),
    .io_storeDataDone_2(loadQ_io_storeDataDone_2),
    .io_storeDataDone_3(loadQ_io_storeDataDone_3),
    .io_storeDataDone_4(loadQ_io_storeDataDone_4),
    .io_storeDataDone_5(loadQ_io_storeDataDone_5),
    .io_storeDataDone_6(loadQ_io_storeDataDone_6),
    .io_storeDataDone_7(loadQ_io_storeDataDone_7),
    .io_storeAddrQueue_0(loadQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(loadQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(loadQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(loadQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(loadQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(loadQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(loadQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(loadQ_io_storeAddrQueue_7),
    .io_storeDataQueue_0(loadQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(loadQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(loadQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(loadQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(loadQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(loadQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(loadQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(loadQ_io_storeDataQueue_7),
    .io_loadAddrDone_0(loadQ_io_loadAddrDone_0),
    .io_loadAddrDone_1(loadQ_io_loadAddrDone_1),
    .io_loadAddrDone_2(loadQ_io_loadAddrDone_2),
    .io_loadAddrDone_3(loadQ_io_loadAddrDone_3),
    .io_loadAddrDone_4(loadQ_io_loadAddrDone_4),
    .io_loadAddrDone_5(loadQ_io_loadAddrDone_5),
    .io_loadAddrDone_6(loadQ_io_loadAddrDone_6),
    .io_loadAddrDone_7(loadQ_io_loadAddrDone_7),
    .io_loadDataDone_0(loadQ_io_loadDataDone_0),
    .io_loadDataDone_1(loadQ_io_loadDataDone_1),
    .io_loadDataDone_2(loadQ_io_loadDataDone_2),
    .io_loadDataDone_3(loadQ_io_loadDataDone_3),
    .io_loadDataDone_4(loadQ_io_loadDataDone_4),
    .io_loadDataDone_5(loadQ_io_loadDataDone_5),
    .io_loadDataDone_6(loadQ_io_loadDataDone_6),
    .io_loadDataDone_7(loadQ_io_loadDataDone_7),
    .io_loadAddrQueue_0(loadQ_io_loadAddrQueue_0),
    .io_loadAddrQueue_1(loadQ_io_loadAddrQueue_1),
    .io_loadAddrQueue_2(loadQ_io_loadAddrQueue_2),
    .io_loadAddrQueue_3(loadQ_io_loadAddrQueue_3),
    .io_loadAddrQueue_4(loadQ_io_loadAddrQueue_4),
    .io_loadAddrQueue_5(loadQ_io_loadAddrQueue_5),
    .io_loadAddrQueue_6(loadQ_io_loadAddrQueue_6),
    .io_loadAddrQueue_7(loadQ_io_loadAddrQueue_7),
    .io_loadAddrEnable_0(loadQ_io_loadAddrEnable_0),
    .io_loadAddrEnable_1(loadQ_io_loadAddrEnable_1),
    .io_addrFromLoadPorts_0(loadQ_io_addrFromLoadPorts_0),
    .io_addrFromLoadPorts_1(loadQ_io_addrFromLoadPorts_1),
    .io_loadPorts_0_ready(loadQ_io_loadPorts_0_ready),
    .io_loadPorts_0_valid(loadQ_io_loadPorts_0_valid),
    .io_loadPorts_0_bits(loadQ_io_loadPorts_0_bits),
    .io_loadPorts_1_ready(loadQ_io_loadPorts_1_ready),
    .io_loadPorts_1_valid(loadQ_io_loadPorts_1_valid),
    .io_loadPorts_1_bits(loadQ_io_loadPorts_1_bits),
    .io_loadDataFromMem(loadQ_io_loadDataFromMem),
    .io_loadAddrToMem(loadQ_io_loadAddrToMem),
    .io_loadEnableToMem(loadQ_io_loadEnableToMem),
    .io_memIsReadyForLoads(loadQ_io_memIsReadyForLoads)
  );
  GROUP_ALLOCATOR_LSQ_A GA ( // @[LSQBRAM.scala 74:18:@12659.4]
    .io_bbLoadOffsets_0(GA_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(GA_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(GA_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(GA_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(GA_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(GA_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(GA_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(GA_io_bbLoadOffsets_7),
    .io_bbLoadPorts_1(GA_io_bbLoadPorts_1),
    .io_bbNumLoads(GA_io_bbNumLoads),
    .io_loadTail(GA_io_loadTail),
    .io_loadHead(GA_io_loadHead),
    .io_loadEmpty(GA_io_loadEmpty),
    .io_bbStoreOffsets_0(GA_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(GA_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(GA_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(GA_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(GA_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(GA_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(GA_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(GA_io_bbStoreOffsets_7),
    .io_bbStorePorts_1(GA_io_bbStorePorts_1),
    .io_bbNumStores(GA_io_bbNumStores),
    .io_storeTail(GA_io_storeTail),
    .io_storeHead(GA_io_storeHead),
    .io_storeEmpty(GA_io_storeEmpty),
    .io_bbStart(GA_io_bbStart),
    .io_bbStartSignals_0(GA_io_bbStartSignals_0),
    .io_readyToPrevious_0(GA_io_readyToPrevious_0),
    .io_loadPortsEnable_0(GA_io_loadPortsEnable_0),
    .io_loadPortsEnable_1(GA_io_loadPortsEnable_1),
    .io_storePortsEnable_0(GA_io_storePortsEnable_0),
    .io_storePortsEnable_1(GA_io_storePortsEnable_1)
  );
  LOAD_PORT_LSQ_A LOAD_PORT_LSQ_A ( // @[LSQBRAM.scala 77:11:@12662.4]
    .clock(LOAD_PORT_LSQ_A_clock),
    .reset(LOAD_PORT_LSQ_A_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_A_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_A_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_A_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_A_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_A_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_A_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_A_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_A_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_A_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_A_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_A_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_A_io_dataFromLoadQueue_bits)
  );
  LOAD_PORT_LSQ_A LOAD_PORT_LSQ_A_1 ( // @[LSQBRAM.scala 77:11:@12665.4]
    .clock(LOAD_PORT_LSQ_A_1_clock),
    .reset(LOAD_PORT_LSQ_A_1_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_A_1_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_A_1_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_A_1_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_A_1_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_A_1_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_A_1_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_A_1_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_A_1_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_A_1_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_A_1_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_A_1_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_A_1_io_dataFromLoadQueue_bits)
  );
  STORE_DATA_PORT_LSQ_A STORE_DATA_PORT_LSQ_A ( // @[LSQBRAM.scala 80:11:@12693.4]
    .clock(STORE_DATA_PORT_LSQ_A_clock),
    .reset(STORE_DATA_PORT_LSQ_A_reset),
    .io_dataFromPrev_ready(STORE_DATA_PORT_LSQ_A_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_DATA_PORT_LSQ_A_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_DATA_PORT_LSQ_A_io_dataFromPrev_bits),
    .io_portEnable(STORE_DATA_PORT_LSQ_A_io_portEnable),
    .io_storeDataEnable(STORE_DATA_PORT_LSQ_A_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_DATA_PORT_LSQ_A_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_A STORE_DATA_PORT_LSQ_A_1 ( // @[LSQBRAM.scala 80:11:@12696.4]
    .clock(STORE_DATA_PORT_LSQ_A_1_clock),
    .reset(STORE_DATA_PORT_LSQ_A_1_reset),
    .io_dataFromPrev_ready(STORE_DATA_PORT_LSQ_A_1_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_DATA_PORT_LSQ_A_1_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_DATA_PORT_LSQ_A_1_io_dataFromPrev_bits),
    .io_portEnable(STORE_DATA_PORT_LSQ_A_1_io_portEnable),
    .io_storeDataEnable(STORE_DATA_PORT_LSQ_A_1_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_DATA_PORT_LSQ_A_1_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_A STORE_ADDR_PORT_LSQ_A ( // @[LSQBRAM.scala 83:11:@12712.4]
    .clock(STORE_ADDR_PORT_LSQ_A_clock),
    .reset(STORE_ADDR_PORT_LSQ_A_reset),
    .io_dataFromPrev_ready(STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_bits),
    .io_portEnable(STORE_ADDR_PORT_LSQ_A_io_portEnable),
    .io_storeDataEnable(STORE_ADDR_PORT_LSQ_A_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_ADDR_PORT_LSQ_A_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_A STORE_ADDR_PORT_LSQ_A_1 ( // @[LSQBRAM.scala 83:11:@12715.4]
    .clock(STORE_ADDR_PORT_LSQ_A_1_clock),
    .reset(STORE_ADDR_PORT_LSQ_A_1_reset),
    .io_dataFromPrev_ready(STORE_ADDR_PORT_LSQ_A_1_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_ADDR_PORT_LSQ_A_1_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_ADDR_PORT_LSQ_A_1_io_dataFromPrev_bits),
    .io_portEnable(STORE_ADDR_PORT_LSQ_A_1_io_portEnable),
    .io_storeDataEnable(STORE_ADDR_PORT_LSQ_A_1_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_ADDR_PORT_LSQ_A_1_io_dataToStoreQueue)
  );
  assign storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 46:24:@12629.4 LSQBRAM.scala 151:14:@12921.4]
  assign loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 52:23:@12635.4 LSQBRAM.scala 119:13:@12835.4]
  assign storeTail = {{5'd0}, storeQ_io_storeTail}; // @[LSQBRAM.scala 44:23:@12627.4 LSQBRAM.scala 149:13:@12919.4]
  assign storeHead = {{5'd0}, storeQ_io_storeHead}; // @[LSQBRAM.scala 45:23:@12628.4 LSQBRAM.scala 150:13:@12920.4]
  assign loadTail = {{5'd0}, loadQ_io_loadTail}; // @[LSQBRAM.scala 50:22:@12633.4 LSQBRAM.scala 117:12:@12833.4]
  assign loadHead = {{5'd0}, loadQ_io_loadHead}; // @[LSQBRAM.scala 51:22:@12634.4 LSQBRAM.scala 118:12:@12834.4]
  assign io_storeDataOut = storeQ_io_storeDataToMem; // @[LSQBRAM.scala 161:19:@12963.4]
  assign io_storeAddrOut = storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 160:19:@12962.4]
  assign io_storeEnable = storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 162:18:@12964.4]
  assign io_loadAddrOut = loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 135:18:@12872.4]
  assign io_loadEnable = loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 136:17:@12873.4]
  assign io_bbReadyToPrevs_0 = GA_io_readyToPrevious_0; // @[LSQBRAM.scala 102:21:@12775.4]
  assign io_rdPortsPrev_0_ready = LOAD_PORT_LSQ_A_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@12968.4]
  assign io_rdPortsPrev_1_ready = LOAD_PORT_LSQ_A_1_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@12980.4]
  assign io_rdPortsNext_0_valid = LOAD_PORT_LSQ_A_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@12971.4]
  assign io_rdPortsNext_0_bits = LOAD_PORT_LSQ_A_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@12970.4]
  assign io_rdPortsNext_1_valid = LOAD_PORT_LSQ_A_1_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@12983.4]
  assign io_rdPortsNext_1_bits = LOAD_PORT_LSQ_A_1_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@12982.4]
  assign io_wrAddrPorts_0_ready = STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_ready; // @[LSQBRAM.scala 182:39:@12998.4]
  assign io_wrAddrPorts_1_ready = STORE_ADDR_PORT_LSQ_A_1_io_dataFromPrev_ready; // @[LSQBRAM.scala 182:39:@13010.4]
  assign io_wrDataPorts_0_ready = STORE_DATA_PORT_LSQ_A_io_dataFromPrev_ready; // @[LSQBRAM.scala 177:36:@12992.4]
  assign io_wrDataPorts_1_ready = STORE_DATA_PORT_LSQ_A_1_io_dataFromPrev_ready; // @[LSQBRAM.scala 177:36:@13004.4]
  assign io_Empty_Valid = storeEmpty & loadEmpty; // @[LSQBRAM.scala 86:18:@12732.4]
  assign storeQ_clock = clock; // @[:@12654.4]
  assign storeQ_reset = reset; // @[:@12655.4]
  assign storeQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 145:21:@12901.4]
  assign storeQ_io_bbStoreOffsets_0 = GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 146:28:@12902.4]
  assign storeQ_io_bbStoreOffsets_1 = GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 146:28:@12903.4]
  assign storeQ_io_bbStoreOffsets_2 = GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 146:28:@12904.4]
  assign storeQ_io_bbStoreOffsets_3 = GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 146:28:@12905.4]
  assign storeQ_io_bbStoreOffsets_4 = GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 146:28:@12906.4]
  assign storeQ_io_bbStoreOffsets_5 = GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 146:28:@12907.4]
  assign storeQ_io_bbStoreOffsets_6 = GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 146:28:@12908.4]
  assign storeQ_io_bbStoreOffsets_7 = GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 146:28:@12909.4]
  assign storeQ_io_bbStorePorts_1 = GA_io_bbStorePorts_1; // @[LSQBRAM.scala 147:26:@12911.4]
  assign storeQ_io_bbNumStores = GA_io_bbNumStores; // @[LSQBRAM.scala 148:25:@12918.4]
  assign storeQ_io_loadTail = loadTail[2:0]; // @[LSQBRAM.scala 139:22:@12874.4]
  assign storeQ_io_loadHead = loadHead[2:0]; // @[LSQBRAM.scala 140:22:@12875.4]
  assign storeQ_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 141:23:@12876.4]
  assign storeQ_io_loadAddressDone_0 = loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 142:29:@12877.4]
  assign storeQ_io_loadAddressDone_1 = loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 142:29:@12878.4]
  assign storeQ_io_loadAddressDone_2 = loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 142:29:@12879.4]
  assign storeQ_io_loadAddressDone_3 = loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 142:29:@12880.4]
  assign storeQ_io_loadAddressDone_4 = loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 142:29:@12881.4]
  assign storeQ_io_loadAddressDone_5 = loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 142:29:@12882.4]
  assign storeQ_io_loadAddressDone_6 = loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 142:29:@12883.4]
  assign storeQ_io_loadAddressDone_7 = loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 142:29:@12884.4]
  assign storeQ_io_loadDataDone_0 = loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 143:26:@12885.4]
  assign storeQ_io_loadDataDone_1 = loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 143:26:@12886.4]
  assign storeQ_io_loadDataDone_2 = loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 143:26:@12887.4]
  assign storeQ_io_loadDataDone_3 = loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 143:26:@12888.4]
  assign storeQ_io_loadDataDone_4 = loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 143:26:@12889.4]
  assign storeQ_io_loadDataDone_5 = loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 143:26:@12890.4]
  assign storeQ_io_loadDataDone_6 = loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 143:26:@12891.4]
  assign storeQ_io_loadDataDone_7 = loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 143:26:@12892.4]
  assign storeQ_io_loadAddressQueue_0 = loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 144:30:@12893.4]
  assign storeQ_io_loadAddressQueue_1 = loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 144:30:@12894.4]
  assign storeQ_io_loadAddressQueue_2 = loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 144:30:@12895.4]
  assign storeQ_io_loadAddressQueue_3 = loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 144:30:@12896.4]
  assign storeQ_io_loadAddressQueue_4 = loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 144:30:@12897.4]
  assign storeQ_io_loadAddressQueue_5 = loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 144:30:@12898.4]
  assign storeQ_io_loadAddressQueue_6 = loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 144:30:@12899.4]
  assign storeQ_io_loadAddressQueue_7 = loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 144:30:@12900.4]
  assign storeQ_io_storeDataEnable_0 = STORE_DATA_PORT_LSQ_A_io_storeDataEnable; // @[LSQBRAM.scala 156:29:@12954.4]
  assign storeQ_io_storeDataEnable_1 = STORE_DATA_PORT_LSQ_A_1_io_storeDataEnable; // @[LSQBRAM.scala 156:29:@12955.4]
  assign storeQ_io_dataFromStorePorts_0 = STORE_DATA_PORT_LSQ_A_io_dataToStoreQueue; // @[LSQBRAM.scala 157:32:@12956.4]
  assign storeQ_io_dataFromStorePorts_1 = STORE_DATA_PORT_LSQ_A_1_io_dataToStoreQueue; // @[LSQBRAM.scala 157:32:@12957.4]
  assign storeQ_io_storeAddrEnable_0 = STORE_ADDR_PORT_LSQ_A_io_storeDataEnable; // @[LSQBRAM.scala 158:29:@12958.4]
  assign storeQ_io_storeAddrEnable_1 = STORE_ADDR_PORT_LSQ_A_1_io_storeDataEnable; // @[LSQBRAM.scala 158:29:@12959.4]
  assign storeQ_io_addressFromStorePorts_0 = STORE_ADDR_PORT_LSQ_A_io_dataToStoreQueue; // @[LSQBRAM.scala 159:35:@12960.4]
  assign storeQ_io_addressFromStorePorts_1 = STORE_ADDR_PORT_LSQ_A_1_io_dataToStoreQueue; // @[LSQBRAM.scala 159:35:@12961.4]
  assign storeQ_io_memIsReadyForStores = io_memIsReadyForStores; // @[LSQBRAM.scala 163:33:@12965.4]
  assign loadQ_clock = clock; // @[:@12657.4]
  assign loadQ_reset = reset; // @[:@12658.4]
  assign loadQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 113:20:@12815.4]
  assign loadQ_io_bbLoadOffsets_0 = GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 114:26:@12816.4]
  assign loadQ_io_bbLoadOffsets_1 = GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 114:26:@12817.4]
  assign loadQ_io_bbLoadOffsets_2 = GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 114:26:@12818.4]
  assign loadQ_io_bbLoadOffsets_3 = GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 114:26:@12819.4]
  assign loadQ_io_bbLoadOffsets_4 = GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 114:26:@12820.4]
  assign loadQ_io_bbLoadOffsets_5 = GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 114:26:@12821.4]
  assign loadQ_io_bbLoadOffsets_6 = GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 114:26:@12822.4]
  assign loadQ_io_bbLoadOffsets_7 = GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 114:26:@12823.4]
  assign loadQ_io_bbLoadPorts_1 = GA_io_bbLoadPorts_1; // @[LSQBRAM.scala 115:24:@12825.4]
  assign loadQ_io_bbNumLoads = GA_io_bbNumLoads; // @[LSQBRAM.scala 116:23:@12832.4]
  assign loadQ_io_storeTail = storeTail[2:0]; // @[LSQBRAM.scala 106:22:@12780.4]
  assign loadQ_io_storeHead = storeHead[2:0]; // @[LSQBRAM.scala 107:22:@12781.4]
  assign loadQ_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 108:23:@12782.4]
  assign loadQ_io_storeAddrDone_0 = storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 109:26:@12783.4]
  assign loadQ_io_storeAddrDone_1 = storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 109:26:@12784.4]
  assign loadQ_io_storeAddrDone_2 = storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 109:26:@12785.4]
  assign loadQ_io_storeAddrDone_3 = storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 109:26:@12786.4]
  assign loadQ_io_storeAddrDone_4 = storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 109:26:@12787.4]
  assign loadQ_io_storeAddrDone_5 = storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 109:26:@12788.4]
  assign loadQ_io_storeAddrDone_6 = storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 109:26:@12789.4]
  assign loadQ_io_storeAddrDone_7 = storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 109:26:@12790.4]
  assign loadQ_io_storeDataDone_0 = storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 110:26:@12791.4]
  assign loadQ_io_storeDataDone_1 = storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 110:26:@12792.4]
  assign loadQ_io_storeDataDone_2 = storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 110:26:@12793.4]
  assign loadQ_io_storeDataDone_3 = storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 110:26:@12794.4]
  assign loadQ_io_storeDataDone_4 = storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 110:26:@12795.4]
  assign loadQ_io_storeDataDone_5 = storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 110:26:@12796.4]
  assign loadQ_io_storeDataDone_6 = storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 110:26:@12797.4]
  assign loadQ_io_storeDataDone_7 = storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 110:26:@12798.4]
  assign loadQ_io_storeAddrQueue_0 = storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 111:27:@12799.4]
  assign loadQ_io_storeAddrQueue_1 = storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 111:27:@12800.4]
  assign loadQ_io_storeAddrQueue_2 = storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 111:27:@12801.4]
  assign loadQ_io_storeAddrQueue_3 = storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 111:27:@12802.4]
  assign loadQ_io_storeAddrQueue_4 = storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 111:27:@12803.4]
  assign loadQ_io_storeAddrQueue_5 = storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 111:27:@12804.4]
  assign loadQ_io_storeAddrQueue_6 = storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 111:27:@12805.4]
  assign loadQ_io_storeAddrQueue_7 = storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 111:27:@12806.4]
  assign loadQ_io_storeDataQueue_0 = storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 112:27:@12807.4]
  assign loadQ_io_storeDataQueue_1 = storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 112:27:@12808.4]
  assign loadQ_io_storeDataQueue_2 = storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 112:27:@12809.4]
  assign loadQ_io_storeDataQueue_3 = storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 112:27:@12810.4]
  assign loadQ_io_storeDataQueue_4 = storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 112:27:@12811.4]
  assign loadQ_io_storeDataQueue_5 = storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 112:27:@12812.4]
  assign loadQ_io_storeDataQueue_6 = storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 112:27:@12813.4]
  assign loadQ_io_storeDataQueue_7 = storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 112:27:@12814.4]
  assign loadQ_io_loadAddrEnable_0 = LOAD_PORT_LSQ_A_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@12864.4]
  assign loadQ_io_loadAddrEnable_1 = LOAD_PORT_LSQ_A_1_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@12869.4]
  assign loadQ_io_addrFromLoadPorts_0 = LOAD_PORT_LSQ_A_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@12863.4]
  assign loadQ_io_addrFromLoadPorts_1 = LOAD_PORT_LSQ_A_1_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@12868.4]
  assign loadQ_io_loadPorts_0_ready = LOAD_PORT_LSQ_A_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@12862.4]
  assign loadQ_io_loadPorts_1_ready = LOAD_PORT_LSQ_A_1_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@12867.4]
  assign loadQ_io_loadDataFromMem = io_loadDataIn; // @[LSQBRAM.scala 133:28:@12870.4]
  assign loadQ_io_memIsReadyForLoads = io_memIsReadyForLoads; // @[LSQBRAM.scala 134:31:@12871.4]
  assign GA_io_loadTail = loadTail[2:0]; // @[LSQBRAM.scala 91:18:@12750.4]
  assign GA_io_loadHead = loadHead[2:0]; // @[LSQBRAM.scala 92:18:@12751.4]
  assign GA_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 93:19:@12752.4]
  assign GA_io_storeTail = storeTail[2:0]; // @[LSQBRAM.scala 97:19:@12770.4]
  assign GA_io_storeHead = storeHead[2:0]; // @[LSQBRAM.scala 98:19:@12771.4]
  assign GA_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 99:20:@12772.4]
  assign GA_io_bbStartSignals_0 = io_bbpValids_0; // @[LSQBRAM.scala 101:24:@12774.4]
  assign LOAD_PORT_LSQ_A_clock = clock; // @[:@12663.4]
  assign LOAD_PORT_LSQ_A_reset = reset; // @[:@12664.4]
  assign LOAD_PORT_LSQ_A_io_addrFromPrev_valid = io_rdPortsPrev_0_valid; // @[LSQBRAM.scala 76:26:@12679.4]
  assign LOAD_PORT_LSQ_A_io_addrFromPrev_bits = io_rdPortsPrev_0_bits; // @[LSQBRAM.scala 76:26:@12678.4]
  assign LOAD_PORT_LSQ_A_io_portEnable = GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 76:26:@12677.4]
  assign LOAD_PORT_LSQ_A_io_dataToNext_ready = io_rdPortsNext_0_ready; // @[LSQBRAM.scala 76:26:@12676.4]
  assign LOAD_PORT_LSQ_A_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 76:26:@12670.4]
  assign LOAD_PORT_LSQ_A_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 76:26:@12669.4]
  assign LOAD_PORT_LSQ_A_1_clock = clock; // @[:@12666.4]
  assign LOAD_PORT_LSQ_A_1_reset = reset; // @[:@12667.4]
  assign LOAD_PORT_LSQ_A_1_io_addrFromPrev_valid = io_rdPortsPrev_1_valid; // @[LSQBRAM.scala 76:26:@12691.4]
  assign LOAD_PORT_LSQ_A_1_io_addrFromPrev_bits = io_rdPortsPrev_1_bits; // @[LSQBRAM.scala 76:26:@12690.4]
  assign LOAD_PORT_LSQ_A_1_io_portEnable = GA_io_loadPortsEnable_1; // @[LSQBRAM.scala 76:26:@12689.4]
  assign LOAD_PORT_LSQ_A_1_io_dataToNext_ready = io_rdPortsNext_1_ready; // @[LSQBRAM.scala 76:26:@12688.4]
  assign LOAD_PORT_LSQ_A_1_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_1_valid; // @[LSQBRAM.scala 76:26:@12682.4]
  assign LOAD_PORT_LSQ_A_1_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_1_bits; // @[LSQBRAM.scala 76:26:@12681.4]
  assign STORE_DATA_PORT_LSQ_A_clock = clock; // @[:@12694.4]
  assign STORE_DATA_PORT_LSQ_A_reset = reset; // @[:@12695.4]
  assign STORE_DATA_PORT_LSQ_A_io_dataFromPrev_valid = io_wrDataPorts_0_valid; // @[LSQBRAM.scala 79:31:@12704.4]
  assign STORE_DATA_PORT_LSQ_A_io_dataFromPrev_bits = io_wrDataPorts_0_bits; // @[LSQBRAM.scala 79:31:@12703.4]
  assign STORE_DATA_PORT_LSQ_A_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 79:31:@12702.4]
  assign STORE_DATA_PORT_LSQ_A_1_clock = clock; // @[:@12697.4]
  assign STORE_DATA_PORT_LSQ_A_1_reset = reset; // @[:@12698.4]
  assign STORE_DATA_PORT_LSQ_A_1_io_dataFromPrev_valid = io_wrDataPorts_1_valid; // @[LSQBRAM.scala 79:31:@12710.4]
  assign STORE_DATA_PORT_LSQ_A_1_io_dataFromPrev_bits = io_wrDataPorts_1_bits; // @[LSQBRAM.scala 79:31:@12709.4]
  assign STORE_DATA_PORT_LSQ_A_1_io_portEnable = GA_io_storePortsEnable_1; // @[LSQBRAM.scala 79:31:@12708.4]
  assign STORE_ADDR_PORT_LSQ_A_clock = clock; // @[:@12713.4]
  assign STORE_ADDR_PORT_LSQ_A_reset = reset; // @[:@12714.4]
  assign STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_valid = io_wrAddrPorts_0_valid; // @[LSQBRAM.scala 82:34:@12723.4]
  assign STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_bits = io_wrAddrPorts_0_bits; // @[LSQBRAM.scala 82:34:@12722.4]
  assign STORE_ADDR_PORT_LSQ_A_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 82:34:@12721.4]
  assign STORE_ADDR_PORT_LSQ_A_1_clock = clock; // @[:@12716.4]
  assign STORE_ADDR_PORT_LSQ_A_1_reset = reset; // @[:@12717.4]
  assign STORE_ADDR_PORT_LSQ_A_1_io_dataFromPrev_valid = io_wrAddrPorts_1_valid; // @[LSQBRAM.scala 82:34:@12729.4]
  assign STORE_ADDR_PORT_LSQ_A_1_io_dataFromPrev_bits = io_wrAddrPorts_1_bits; // @[LSQBRAM.scala 82:34:@12728.4]
  assign STORE_ADDR_PORT_LSQ_A_1_io_portEnable = GA_io_storePortsEnable_1; // @[LSQBRAM.scala 82:34:@12727.4]
endmodule
